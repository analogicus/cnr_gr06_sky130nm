magic
tech sky130B
magscale 1 2
timestamp 1713382108
<< checkpaint >>
rect -1313 6192 1799 6245
rect -1313 6139 2338 6192
rect -1313 6086 2877 6139
rect -1313 6033 3416 6086
rect -1313 5980 3955 6033
rect -1313 5927 4494 5980
rect -1313 5874 5033 5927
rect -1313 5662 5572 5874
rect -1313 -713 7728 5662
rect -1260 -978 7728 -713
rect -1260 -3660 1460 -978
rect 1921 -1031 7728 -978
rect 2460 -1084 7728 -1031
rect 4616 -1296 7728 -1084
<< error_s >>
rect 468 4915 503 4949
rect 469 4896 503 4915
rect 488 583 503 4896
rect 522 4862 557 4896
rect 1007 4862 1042 4896
rect 522 583 556 4862
rect 1008 4843 1042 4862
rect 522 549 537 583
rect 1027 530 1042 4843
rect 1061 4809 1096 4843
rect 1546 4809 1581 4843
rect 1061 530 1095 4809
rect 1547 4790 1581 4809
rect 1061 496 1076 530
rect 1566 477 1581 4790
rect 1600 4756 1635 4790
rect 2085 4756 2120 4790
rect 1600 477 1634 4756
rect 2086 4737 2120 4756
rect 1600 443 1615 477
rect 2105 424 2120 4737
rect 2139 4703 2174 4737
rect 2624 4703 2659 4737
rect 2139 424 2173 4703
rect 2625 4684 2659 4703
rect 2139 390 2154 424
rect 2644 371 2659 4684
rect 2678 4650 2713 4684
rect 3163 4650 3198 4684
rect 2678 371 2712 4650
rect 3164 4631 3198 4650
rect 2678 337 2693 371
rect 3183 318 3198 4631
rect 3217 4597 3252 4631
rect 3702 4597 3737 4631
rect 3217 318 3251 4597
rect 3703 4578 3737 4597
rect 3217 284 3232 318
rect 3722 265 3737 4578
rect 3756 4544 3791 4578
rect 3756 265 3790 4544
rect 4242 2543 4276 2561
rect 4242 2507 4312 2543
rect 4259 2473 4330 2507
rect 4780 2473 4815 2507
rect 3756 231 3771 265
rect 4259 212 4329 2473
rect 4781 2454 4815 2473
rect 4259 176 4312 212
rect 4800 159 4815 2454
rect 4834 2420 4869 2454
rect 5319 2420 5354 2454
rect 5912 2437 5946 2455
rect 4834 159 4868 2420
rect 5320 2401 5354 2420
rect 4834 125 4849 159
rect 5339 106 5354 2401
rect 5373 2367 5408 2401
rect 5373 106 5407 2367
rect 5373 72 5388 106
rect 5876 53 5946 2437
rect 6398 2331 6432 2349
rect 6398 2295 6468 2331
rect 6415 2261 6486 2295
rect 6936 2261 6971 2295
rect 5876 17 5929 53
rect 6415 0 6485 2261
rect 6937 2242 6971 2261
rect 6415 -36 6468 0
rect 6956 -53 6971 2242
rect 6990 2208 7025 2242
rect 6990 -53 7024 2208
rect 6990 -87 7005 -53
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
use sky130_fd_pr__pfet_01v8_6HSZAW  XM1
timestamp 0
transform 1 0 243 0 1 2766
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM2
timestamp 0
transform 1 0 782 0 1 2713
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM3
timestamp 0
transform 1 0 1321 0 1 2660
box -296 -2219 296 2219
use sky130_fd_pr__nfet_01v8_6WXQK8  XM4
timestamp 0
transform 1 0 7250 0 1 1068
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_6HSZAW  XM5
timestamp 0
transform 1 0 1860 0 1 2607
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM6
timestamp 0
transform 1 0 2399 0 1 2554
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM7
timestamp 0
transform 1 0 2938 0 1 2501
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM8
timestamp 0
transform 1 0 3477 0 1 2448
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM9
timestamp 0
transform 1 0 4016 0 1 2395
box -296 -2219 296 2219
use sky130_fd_pr__nfet_01v8_6WXQK8  XM10
timestamp 0
transform 1 0 4555 0 1 1333
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM11
timestamp 0
transform 1 0 5094 0 1 1280
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM12
timestamp 0
transform 1 0 5633 0 1 1227
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_6HSZAW  XM13
timestamp 0
transform 1 0 6172 0 1 2183
box -296 -2219 296 2219
use sky130_fd_pr__nfet_01v8_6WXQK8  XM14
timestamp 0
transform 1 0 6711 0 1 1121
box -296 -1210 296 1210
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD_1V8
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Clk
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vocn
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vocp
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 Vref_c
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Vin_c
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 VSS
port 6 nsew
<< end >>
