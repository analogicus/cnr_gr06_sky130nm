** sch_path: /home/alvaros/aicex/ip/cnr_gr06_sky130nm/design/CNR_GR06_SKY130NM/CNR_GR06_test.sch
**.subckt CNR_GR06_test VDD_1V8 VSS Vn Vp
*.ipin VDD_1V8
*.ipin VSS
*.opin Vn
*.opin Vp
x3 net10 net1 VDD_1V8 VDD_1V8 SUNTR_PCHLCM
x4 net2 net1 VDD_1V8 VDD_1V8 SUNTR_PCHLCM
x5 net4 net1 VDD_1V8 VDD_1V8 SUNTR_PCHLCM
x6 net11 net1 VDD_1V8 VDD_1V8 SUNTR_PCHLCM
x7 Vn net1 VDD_1V8 VDD_1V8 SUNTR_PCHLCM
x8 net6 net7 VDD_1V8 VDD_1V8 SUNTR_PCHLCM
x9 net7 net7 net6 VDD_1V8 SUNTR_PCHLCM
x10 net9 Vp net7 VDD_1V8 SUNTR_PCHLCM
x11 Vp Vp net6 VDD_1V8 SUNTR_PCHLCM
x12 Vp net8 VSS VSS SUNTR_NCHLCM
x13 net9 net8 VSS VSS SUNTR_NCHLCM
x14 Vn Vn net5 VSS SUNTR_NCHLCM
x15 net12 net12 net5 VSS SUNTR_NCHLCM
x16 net5 net12 VSS VSS SUNTR_NCHLCM
x17 net11 Vn net12 VSS SUNTR_NCHLCM
x18 net4 net4 VSS VSS SUNTR_NCHLCM
x19 net3 net4 VSS VSS SUNTR_NCHLCM
x20 net2 net10 net13 VSS SUNTR_NCHLCM
x21 net10 net10 VSS VSS SUNTR_NCHLCM
**.ends

* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_PCHLCM.sym # of pins=4
** sym_path: /home/alvaros/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHLCM.sym
** sch_path: /home/alvaros/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHLCM.sch
.subckt SUNTR_PCHLCM D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM0 N0 G S B SUNTR_PCHL
XM7 D G N0 B SUNTR_PCHL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NCHLCM.sym # of pins=4
** sym_path: /home/alvaros/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHLCM.sym
** sch_path: /home/alvaros/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHLCM.sch
.subckt SUNTR_NCHLCM D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM0 N0 G S B SUNTR_NCHL
XM1 N1 G N0 B SUNTR_NCHL
XM2 N2 G N1 B SUNTR_NCHL
XM3 N3 G N2 B SUNTR_NCHL
XM6 N6 G N3 B SUNTR_NCHL
XM7 N7 G N6 B SUNTR_NCHL
XM8 D G N7 B SUNTR_NCHL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_PCHL.sym # of pins=4
** sym_path: /home/alvaros/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHL.sym
** sch_path: /home/alvaros/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHL.sch
.subckt SUNTR_PCHL D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.36 W=1.08 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NCHL.sym # of pins=4
** sym_path: /home/alvaros/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHL.sym
** sch_path: /home/alvaros/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHL.sch
.subckt SUNTR_NCHL D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.36 W=1.08 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
