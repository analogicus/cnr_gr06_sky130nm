magic
tech sky130B
magscale 1 2
timestamp 1713382108
<< checkpaint >>
rect 5694 5503 8806 5556
rect 5694 5450 9345 5503
rect 5694 5397 9884 5450
rect 5694 5344 10423 5397
rect 5694 5291 10962 5344
rect 5694 5238 11501 5291
rect 5694 5185 12040 5238
rect 5694 5132 12579 5185
rect 5694 5079 13118 5132
rect 5694 5026 13657 5079
rect 5694 4973 14196 5026
rect 5694 4920 14735 4973
rect 5694 4867 15274 4920
rect -1260 -2460 1460 1460
rect 5694 -1402 15813 4867
rect 6233 -1455 15813 -1402
rect 6772 -1508 15813 -1455
rect 7311 -1561 15813 -1508
rect 7850 -1614 15813 -1561
rect 8389 -1667 15813 -1614
rect 8928 -1720 15813 -1667
rect 9467 -1773 15813 -1720
rect 10006 -1826 15813 -1773
rect 10545 -1879 15813 -1826
rect 11084 -1932 15813 -1879
rect 11623 -1985 15813 -1932
rect 12162 -2038 15813 -1985
rect 12701 -2091 15813 -2038
<< error_s >>
rect 7475 4226 7510 4260
rect 7476 4207 7510 4226
rect 468 2897 503 2931
rect 469 2878 503 2897
rect 488 583 503 2878
rect 522 2844 557 2878
rect 1007 2844 1042 2878
rect 522 583 556 2844
rect 1008 2825 1042 2844
rect 522 549 537 583
rect 1027 530 1042 2825
rect 1061 2791 1096 2825
rect 1546 2791 1581 2825
rect 1061 530 1095 2791
rect 1547 2772 1581 2791
rect 1061 496 1076 530
rect 1566 477 1581 2772
rect 1600 2738 1635 2772
rect 2085 2738 2120 2772
rect 1600 477 1634 2738
rect 2086 2719 2120 2738
rect 1600 443 1615 477
rect 2105 424 2120 2719
rect 2139 2685 2174 2719
rect 2624 2685 2659 2719
rect 2139 424 2173 2685
rect 2625 2666 2659 2685
rect 2139 390 2154 424
rect 2644 371 2659 2666
rect 2678 2632 2713 2666
rect 3163 2632 3198 2666
rect 2678 371 2712 2632
rect 3164 2613 3198 2632
rect 2678 337 2693 371
rect 3183 318 3198 2613
rect 3217 2579 3252 2613
rect 3702 2579 3737 2613
rect 3217 318 3251 2579
rect 3703 2560 3737 2579
rect 3217 284 3232 318
rect 3722 265 3737 2560
rect 3756 2526 3791 2560
rect 4241 2526 4276 2560
rect 3756 265 3790 2526
rect 4242 2507 4276 2526
rect 3756 231 3771 265
rect 4261 212 4276 2507
rect 4295 2473 4330 2507
rect 4780 2473 4815 2507
rect 4295 212 4329 2473
rect 4781 2454 4815 2473
rect 4295 178 4310 212
rect 4800 159 4815 2454
rect 4834 2420 4869 2454
rect 5319 2420 5354 2454
rect 4834 159 4868 2420
rect 5320 2401 5354 2420
rect 4834 125 4849 159
rect 5339 106 5354 2401
rect 5373 2367 5408 2401
rect 5858 2367 5893 2401
rect 5373 106 5407 2367
rect 5859 2348 5893 2367
rect 5373 72 5388 106
rect 5878 53 5893 2348
rect 5912 2314 5947 2348
rect 6397 2314 6432 2348
rect 6990 2331 7024 2349
rect 5912 53 5946 2314
rect 6398 2295 6432 2314
rect 5912 19 5927 53
rect 6417 0 6432 2295
rect 6451 2261 6486 2295
rect 6451 0 6485 2261
rect 6451 -34 6466 0
rect 6954 -53 7024 2331
rect 6954 -89 7007 -53
rect 7495 -106 7510 4207
rect 7529 4173 7564 4207
rect 8014 4173 8049 4207
rect 7529 -106 7563 4173
rect 8015 4154 8049 4173
rect 7529 -140 7544 -106
rect 8034 -159 8049 4154
rect 8068 4120 8103 4154
rect 8553 4120 8588 4154
rect 8068 -159 8102 4120
rect 8554 4101 8588 4120
rect 8068 -193 8083 -159
rect 8573 -212 8588 4101
rect 8607 4067 8642 4101
rect 9092 4067 9127 4101
rect 8607 -212 8641 4067
rect 9093 4048 9127 4067
rect 8607 -246 8622 -212
rect 9112 -265 9127 4048
rect 9146 4014 9181 4048
rect 9631 4014 9666 4048
rect 9146 -265 9180 4014
rect 9632 3995 9666 4014
rect 9146 -299 9161 -265
rect 9651 -318 9666 3995
rect 9685 3961 9720 3995
rect 10170 3961 10205 3995
rect 9685 -318 9719 3961
rect 10171 3942 10205 3961
rect 9685 -352 9700 -318
rect 10190 -371 10205 3942
rect 10224 3908 10259 3942
rect 10709 3908 10744 3942
rect 10224 -371 10258 3908
rect 10710 3889 10744 3908
rect 10224 -405 10239 -371
rect 10729 -424 10744 3889
rect 10763 3855 10798 3889
rect 11248 3855 11283 3889
rect 10763 -424 10797 3855
rect 11249 3836 11283 3855
rect 10763 -458 10778 -424
rect 11268 -477 11283 3836
rect 11302 3802 11337 3836
rect 11787 3802 11822 3836
rect 11302 -477 11336 3802
rect 11788 3783 11822 3802
rect 11302 -511 11317 -477
rect 11807 -530 11822 3783
rect 11841 3749 11876 3783
rect 12326 3749 12361 3783
rect 11841 -530 11875 3749
rect 12327 3730 12361 3749
rect 11841 -564 11856 -530
rect 12346 -583 12361 3730
rect 12380 3696 12415 3730
rect 12865 3696 12900 3730
rect 12380 -583 12414 3696
rect 12866 3677 12900 3696
rect 12380 -617 12395 -583
rect 12885 -636 12900 3677
rect 12919 3643 12954 3677
rect 13404 3643 13439 3677
rect 12919 -636 12953 3643
rect 13405 3624 13439 3643
rect 12919 -670 12934 -636
rect 13424 -689 13439 3624
rect 13458 3590 13493 3624
rect 13943 3590 13978 3624
rect 13458 -689 13492 3590
rect 13944 3571 13978 3590
rect 13458 -723 13473 -689
rect 13963 -742 13978 3571
rect 13997 3537 14032 3571
rect 13997 -742 14031 3537
rect 13997 -776 14012 -742
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__nfet_01v8_6WXQK8  XM1
timestamp 0
transform 1 0 243 0 1 1757
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM2
timestamp 0
transform 1 0 782 0 1 1704
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM3
timestamp 0
transform 1 0 1321 0 1 1651
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_6HSZAW  XM4
timestamp 0
transform 1 0 7250 0 1 2077
box -296 -2219 296 2219
use sky130_fd_pr__nfet_01v8_6WXQK8  XM5
timestamp 0
transform 1 0 1860 0 1 1598
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM6
timestamp 0
transform 1 0 2399 0 1 1545
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM7
timestamp 0
transform 1 0 2938 0 1 1492
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM8
timestamp 0
transform 1 0 3477 0 1 1439
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM9
timestamp 0
transform 1 0 4016 0 1 1386
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM10
timestamp 0
transform 1 0 4555 0 1 1333
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM11
timestamp 0
transform 1 0 5094 0 1 1280
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM12
timestamp 0
transform 1 0 5633 0 1 1227
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM13
timestamp 0
transform 1 0 6172 0 1 1174
box -296 -1210 296 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  XM14
timestamp 0
transform 1 0 6711 0 1 1121
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_6HSZAW  XM15
timestamp 0
transform 1 0 7789 0 1 2024
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM16
timestamp 0
transform 1 0 8328 0 1 1971
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM17
timestamp 0
transform 1 0 8867 0 1 1918
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM18
timestamp 0
transform 1 0 9406 0 1 1865
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM19
timestamp 0
transform 1 0 9945 0 1 1812
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM20
timestamp 0
transform 1 0 10484 0 1 1759
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM21
timestamp 0
transform 1 0 11023 0 1 1706
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM22
timestamp 0
transform 1 0 11562 0 1 1653
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM23
timestamp 0
transform 1 0 12101 0 1 1600
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM24
timestamp 0
transform 1 0 12640 0 1 1547
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM25
timestamp 0
transform 1 0 13179 0 1 1494
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM26
timestamp 0
transform 1 0 13718 0 1 1441
box -296 -2219 296 2219
use sky130_fd_pr__pfet_01v8_6HSZAW  XM27
timestamp 0
transform 1 0 14257 0 1 1388
box -296 -2219 296 2219
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD_1V8
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vn
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vp
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VSS
port 3 nsew
<< end >>
