*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR06_main_lpe.spi
#else
.include ../../../work/xsch/CNR_GR06_main.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 100p

.param t_start = 0.5u
.param t_start_del = {t_start + TRF}

*- 8 MHz clock frequency
.param PERIOD_CLK = 500n

*- 25% duty-cycle clock
.param PW_CLK = PERIOD_CLK/2

*- Supply, vdda is set in includes
.param AVDD = {vdda}
*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0  dc 0
VDD  VDD_1V8 0 dc 1.2
Vdref Vdref 0 dc 0.8

*VT2 VT2 0 dc 0.4
*VT1 VT1 0 dc 0.45

VT1 VT1 0 dc 0 pulse -0.2 0.2 {t_start} {TRF} {TRF} {10000n/2} {10000n}
VT2 VT2 0 dc 0 pulse -0.2 0.2 {t_start+5000n} {TRF} {TRF} {10000n/2} {10000n}

*VT2  VT2 0 SIN(0 0.150 50000 0 0 180)
*VT1  VT1 0 SIN(0 0.150 50000 0 0)

VBP VBP 0 dc 0.144
VBN VBN 0 dc 1.08

VCLK Clk 0 dc 0 pulse 0 1.2 {t_start} {TRF} {TRF} {PW_CLK} {PERIOD_CLK}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save ${VPORTS}
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

tran 0.1u 30u 0.5u
write
quit

.endc

.end
