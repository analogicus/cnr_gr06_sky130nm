*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR06_main_lpe.spi
#else
.include ../../../work/xsch/CNR_GR06_main.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 100p
.param t_start = 0.5u
.param t_start_del = {t_start + TRF}
.param PERIOD_CLK = 500n
.param PW_CLK = PERIOD_CLK/2
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0  dc 0
VDD  VDD_1V8 0 dc 1.2
Vdref Vdref 0 dc 1.2

VT2  VT2 0 SIN(0 0.25 10000 0 0 180)
VT1  VT1 0 SIN(0 0.25 10000 0 0)

VBP VBP 0 dc 0.08
VBN VBN 0 dc 1.12

VCLK Clk 0 dc 0 pulse 0 1.2 {t_start} {TRF} {TRF} {PW_CLK} {PERIOD_CLK}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
#ifdef Debug
.save all
#else
.save ${VPORTS}
#endif

*----------------------------------------------------------------
* NGSPICE control for illustrative purposes (Not actual Monte Carlo)
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

* Just a demonstration loop - not actual Monte Carlo in ngspice context
let runs = 1000
do i = 1, runs
    * Here you would inject randomized parameters externally
    run
    set filetype=ascii
    * This would ideally output to a different file each time
    write "output_data_${i}.txt" V(Voc)
end

.quit
.endc

.end

