magic
tech sky130B
magscale 1 2
timestamp 1713382353
<< error_s >>
rect 147 1045 211 1051
rect 147 1011 159 1045
rect 147 1005 211 1011
rect 147 719 211 725
rect 147 685 159 719
rect 147 679 211 685
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__nfet_01v8_DLP4BZ  XM1
timestamp 1713382353
transform 1 0 179 0 1 865
box -232 -318 232 318
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 D
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 G
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 S
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 B
port 3 nsew
<< end >>
