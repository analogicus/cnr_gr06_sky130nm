magic
tech sky130B
magscale 1 2
timestamp 1713381689
<< checkpaint >>
rect -1313 -1366366 1799 -1366313
rect -1313 -1366419 2338 -1366366
rect -1313 -1366472 2877 -1366419
rect -1313 -1366525 3416 -1366472
rect -1313 -1366578 3955 -1366525
rect -1313 -1366631 4494 -1366578
rect -1313 -1366684 5033 -1366631
rect -1313 -1369353 5572 -1366684
rect -774 -1369406 5572 -1369353
rect -235 -1369459 5572 -1369406
rect 304 -1369512 5572 -1369459
rect 843 -1369565 5572 -1369512
rect 1382 -1369618 5572 -1369565
rect 1921 -1369671 5572 -1369618
rect 2460 -1369724 5572 -1369671
<< error_p >>
rect 40060 -1357631 40095 -1357597
rect 40061 -1357650 40095 -1357631
rect 40080 -1357905 40095 -1357650
rect 40114 -1357684 40149 -1357650
rect 40599 -1357684 40634 -1357650
rect 40114 -1357905 40148 -1357684
rect 40600 -1357703 40634 -1357684
rect 40619 -1357905 40634 -1357703
rect 40653 -1357737 40688 -1357703
rect 41138 -1357737 41173 -1357703
rect 40653 -1357905 40687 -1357737
rect 41139 -1357756 41173 -1357737
rect 41158 -1357905 41173 -1357756
rect 41192 -1357790 41227 -1357756
rect 41677 -1357790 41712 -1357756
rect 41192 -1357905 41226 -1357790
rect 41678 -1357809 41712 -1357790
rect 41697 -1357905 41712 -1357809
rect 41731 -1357843 41766 -1357809
rect 41731 -1357905 41765 -1357843
rect 1546 -1360431 1581 -1360397
rect 1547 -1360450 1581 -1360431
rect 469 -1362326 503 -1362308
rect 1061 -1362326 1095 -1362308
rect 469 -1362362 539 -1362326
rect 486 -1362396 557 -1362362
rect 486 -1364657 556 -1362396
rect 486 -1364693 539 -1364657
rect 1025 -1364710 1095 -1362326
rect 1025 -1364746 1078 -1364710
rect 1566 -1364763 1581 -1360450
rect 1600 -1360484 1635 -1360450
rect 2085 -1360484 2120 -1360450
rect 1600 -1364763 1634 -1360484
rect 2086 -1360503 2120 -1360484
rect 1600 -1364797 1615 -1364763
rect 2105 -1364816 2120 -1360503
rect 2139 -1360537 2174 -1360503
rect 2624 -1360537 2659 -1360503
rect 2139 -1364816 2173 -1360537
rect 2625 -1360556 2659 -1360537
rect 2139 -1364850 2154 -1364816
rect 2644 -1364869 2659 -1360556
rect 2678 -1360590 2713 -1360556
rect 3163 -1360590 3198 -1360556
rect 2678 -1364869 2712 -1360590
rect 3164 -1360609 3198 -1360590
rect 2678 -1364903 2693 -1364869
rect 3183 -1364922 3198 -1360609
rect 3217 -1360643 3252 -1360609
rect 3217 -1364922 3251 -1360643
rect 3703 -1362644 3737 -1362626
rect 3703 -1362680 3773 -1362644
rect 3720 -1362714 3791 -1362680
rect 4241 -1362714 4276 -1362680
rect 3217 -1364956 3232 -1364922
rect 3720 -1364975 3790 -1362714
rect 4242 -1362733 4276 -1362714
rect 3720 -1365011 3773 -1364975
rect 4261 -1365028 4276 -1362733
rect 4295 -1362767 4330 -1362733
rect 4780 -1362767 4815 -1362733
rect 4295 -1365028 4329 -1362767
rect 4781 -1362786 4815 -1362767
rect 4295 -1365062 4310 -1365028
rect 4800 -1365081 4815 -1362786
rect 4834 -1362820 4869 -1362786
rect 5319 -1362820 5354 -1362786
rect 4834 -1365081 4868 -1362820
rect 5320 -1362839 5354 -1362820
rect 4834 -1365115 4849 -1365081
rect 5339 -1365134 5354 -1362839
rect 5373 -1362873 5408 -1362839
rect 5858 -1362873 5893 -1362839
rect 5373 -1365134 5407 -1362873
rect 5859 -1362892 5893 -1362873
rect 5373 -1365168 5388 -1365134
rect 5878 -1365187 5893 -1362892
rect 5912 -1362926 5947 -1362892
rect 6397 -1362926 6432 -1362892
rect 5912 -1365187 5946 -1362926
rect 6398 -1362945 6432 -1362926
rect 5912 -1365221 5927 -1365187
rect 6417 -1365240 6432 -1362945
rect 6451 -1362979 6486 -1362945
rect 6936 -1362979 6971 -1362945
rect 6451 -1365240 6485 -1362979
rect 6937 -1362998 6971 -1362979
rect 6451 -1365274 6466 -1365240
rect 6956 -1365293 6971 -1362998
rect 6990 -1363032 7025 -1362998
rect 6990 -1365293 7024 -1363032
rect 6990 -1365327 7005 -1365293
<< error_s >>
rect 6371 -163840 6372 -157759
rect 12743 -423080 12744 -416999
rect 19115 -587520 19116 -581439
rect 25487 -846720 25488 -840679
rect 31859 -1106000 31860 -1099919
rect 38410 -1361840 38432 -1361640
rect 38438 -1361840 38460 -1361640
rect 38611 -1361840 38638 -1361640
rect 38639 -1361840 38666 -1361640
rect 38812 -1361840 38839 -1361640
rect 38840 -1361840 38867 -1361640
rect 39013 -1361840 39040 -1361640
rect 39041 -1361840 39068 -1361640
rect 39219 -1361840 39241 -1361640
rect 39247 -1361840 39269 -1361640
rect 39425 -1361840 39447 -1361640
rect 39453 -1361840 39475 -1361640
rect 39626 -1361840 39653 -1361640
rect 39654 -1361840 39681 -1361640
rect 39827 -1361840 39854 -1361640
rect 39855 -1361840 39882 -1361640
rect 40033 -1361840 40055 -1361640
rect 40061 -1361840 40083 -1361640
rect 40239 -1361840 40261 -1361640
rect 40267 -1361840 40289 -1361640
rect 40445 -1361840 40467 -1361640
rect 40473 -1361840 40495 -1361640
rect 40646 -1361840 40673 -1361640
rect 40674 -1361840 40701 -1361640
rect 40852 -1361840 40874 -1361640
rect 40880 -1361840 40902 -1361640
rect 41053 -1361840 41080 -1361640
rect 41081 -1361840 41108 -1361640
rect 41259 -1361840 41281 -1361640
rect 41287 -1361840 41309 -1361640
rect 41460 -1361840 41487 -1361640
rect 41488 -1361840 41515 -1361640
rect 41666 -1361840 41688 -1361640
rect 41694 -1361840 41716 -1361640
rect 41867 -1361840 41894 -1361640
rect 41895 -1361840 41922 -1361640
rect 42073 -1361840 42095 -1361640
rect 42101 -1361840 42123 -1361640
rect 42274 -1361840 42301 -1361640
rect 42302 -1361840 42329 -1361640
rect 42480 -1361840 42502 -1361640
rect 42508 -1361840 42530 -1361640
rect 42686 -1361840 42708 -1361640
rect 42714 -1361840 42736 -1361640
rect 42887 -1361840 42914 -1361640
rect 42915 -1361840 42942 -1361640
rect 43088 -1361840 43115 -1361640
rect 43116 -1361840 43143 -1361640
rect 43294 -1361840 43316 -1361640
rect 43322 -1361840 43344 -1361640
rect 43495 -1361840 43522 -1361640
rect 43523 -1361840 43550 -1361640
rect 43701 -1361840 43723 -1361640
rect 43729 -1361840 43751 -1361640
rect 43902 -1361840 43929 -1361640
rect 43930 -1361840 43957 -1361640
rect 44108 -1361840 44130 -1361640
rect 44136 -1361840 44158 -1361640
rect 44309 -1361840 44336 -1361640
rect 44337 -1361840 44364 -1361640
rect 44515 -1361840 44537 -1361640
rect 44543 -1361840 44565 -1361640
rect 44716 -1361840 44743 -1361640
rect 44744 -1361840 44771 -1361640
rect 44922 -1361840 44944 -1361640
rect 44950 -1361840 44972 -1361640
rect 45123 -1361840 45150 -1361640
rect 45151 -1361840 45178 -1361640
rect 45329 -1361840 45351 -1361640
rect 45357 -1361840 45379 -1361640
rect 45530 -1361840 45557 -1361640
rect 45558 -1361840 45585 -1361640
rect 45736 -1361840 45758 -1361640
rect 45764 -1361840 45786 -1361640
rect 45937 -1361840 45964 -1361640
rect 45965 -1361840 45992 -1361640
rect 46143 -1361840 46165 -1361640
rect 46171 -1361840 46193 -1361640
rect 46344 -1361840 46371 -1361640
rect 46372 -1361840 46399 -1361640
rect 46550 -1361840 46572 -1361640
rect 46578 -1361840 46600 -1361640
rect 46751 -1361840 46778 -1361640
rect 46779 -1361840 46806 -1361640
rect 46957 -1361840 46979 -1361640
rect 46985 -1361840 47007 -1361640
rect 47158 -1361840 47185 -1361640
rect 47186 -1361840 47213 -1361640
rect 47364 -1361840 47386 -1361640
rect 47392 -1361840 47414 -1361640
rect 47565 -1361840 47592 -1361640
rect 47593 -1361840 47620 -1361640
rect 47771 -1361840 47793 -1361640
rect 47799 -1361840 47821 -1361640
rect 47972 -1361840 47999 -1361640
rect 48000 -1361840 48027 -1361640
rect 48178 -1361840 48200 -1361640
rect 48206 -1361840 48228 -1361640
rect 48379 -1361840 48406 -1361640
rect 48407 -1361840 48434 -1361640
rect 48585 -1361840 48607 -1361640
rect 48613 -1361840 48635 -1361640
rect 48786 -1361840 48813 -1361640
rect 48814 -1361840 48841 -1361640
rect 48992 -1361840 49014 -1361640
rect 49020 -1361840 49042 -1361640
rect 49193 -1361840 49220 -1361640
rect 49221 -1361840 49248 -1361640
rect 49399 -1361840 49421 -1361640
rect 49427 -1361840 49449 -1361640
rect 49600 -1361840 49627 -1361640
rect 49628 -1361840 49655 -1361640
rect 49806 -1361840 49828 -1361640
rect 49834 -1361840 49856 -1361640
rect 50007 -1361840 50034 -1361640
rect 50035 -1361840 50062 -1361640
rect 50213 -1361840 50235 -1361640
rect 50241 -1361840 50263 -1361640
rect 50414 -1361840 50441 -1361640
rect 50442 -1361840 50469 -1361640
rect 50620 -1361840 50642 -1361640
rect 50648 -1361840 50670 -1361640
rect 50821 -1361840 50848 -1361640
rect 50849 -1361840 50876 -1361640
rect 51027 -1361840 51049 -1361640
rect 51055 -1361840 51077 -1361640
rect 51228 -1361840 51255 -1361640
rect 51256 -1361840 51283 -1361640
rect 51434 -1361840 51456 -1361640
rect 51462 -1361840 51484 -1361640
rect 51635 -1361840 51662 -1361640
rect 51663 -1361840 51690 -1361640
rect 51841 -1361840 51863 -1361640
rect 51869 -1361840 51891 -1361640
rect 52042 -1361840 52069 -1361640
rect 52070 -1361840 52097 -1361640
rect 52248 -1361840 52270 -1361640
rect 52276 -1361840 52298 -1361640
rect 52449 -1361840 52476 -1361640
rect 52477 -1361840 52504 -1361640
rect 52655 -1361840 52677 -1361640
rect 52683 -1361840 52705 -1361640
rect 52856 -1361840 52883 -1361640
rect 52884 -1361840 52911 -1361640
rect 53062 -1361840 53084 -1361640
rect 53090 -1361840 53112 -1361640
rect 53263 -1361840 53290 -1361640
rect 53291 -1361840 53318 -1361640
rect 53469 -1361840 53491 -1361640
rect 53497 -1361840 53519 -1361640
rect 53670 -1361840 53697 -1361640
rect 53698 -1361840 53725 -1361640
rect 53876 -1361840 53898 -1361640
rect 53904 -1361840 53926 -1361640
rect 38410 -1362240 38432 -1362040
rect 38438 -1362240 38460 -1362040
rect 38611 -1362240 38638 -1362040
rect 38639 -1362240 38666 -1362040
rect 38812 -1362240 38839 -1362040
rect 38840 -1362240 38867 -1362040
rect 39013 -1362240 39040 -1362040
rect 39041 -1362240 39068 -1362040
rect 39219 -1362240 39241 -1362040
rect 39247 -1362240 39269 -1362040
rect 39425 -1362240 39447 -1362040
rect 39453 -1362240 39475 -1362040
rect 39626 -1362240 39653 -1362040
rect 39654 -1362240 39681 -1362040
rect 39827 -1362240 39854 -1362040
rect 39855 -1362240 39882 -1362040
rect 40033 -1362240 40055 -1362040
rect 40061 -1362240 40083 -1362040
rect 40239 -1362240 40261 -1362040
rect 40267 -1362240 40289 -1362040
rect 40445 -1362240 40467 -1362040
rect 40473 -1362240 40495 -1362040
rect 40646 -1362240 40673 -1362040
rect 40674 -1362240 40701 -1362040
rect 40852 -1362240 40874 -1362040
rect 40880 -1362240 40902 -1362040
rect 41053 -1362240 41080 -1362040
rect 41081 -1362240 41108 -1362040
rect 41259 -1362240 41281 -1362040
rect 41287 -1362240 41309 -1362040
rect 41460 -1362240 41487 -1362040
rect 41488 -1362240 41515 -1362040
rect 41666 -1362240 41688 -1362040
rect 41694 -1362240 41716 -1362040
rect 41867 -1362240 41894 -1362040
rect 41895 -1362240 41922 -1362040
rect 42073 -1362240 42095 -1362040
rect 42101 -1362240 42123 -1362040
rect 42274 -1362240 42301 -1362040
rect 42302 -1362240 42329 -1362040
rect 42480 -1362240 42502 -1362040
rect 42508 -1362240 42530 -1362040
rect 42686 -1362240 42708 -1362040
rect 42714 -1362240 42736 -1362040
rect 42887 -1362240 42914 -1362040
rect 42915 -1362240 42942 -1362040
rect 43088 -1362240 43115 -1362040
rect 43116 -1362240 43143 -1362040
rect 43294 -1362240 43316 -1362040
rect 43322 -1362240 43344 -1362040
rect 43495 -1362240 43522 -1362040
rect 43523 -1362240 43550 -1362040
rect 43701 -1362240 43723 -1362040
rect 43729 -1362240 43751 -1362040
rect 43902 -1362240 43929 -1362040
rect 43930 -1362240 43957 -1362040
rect 44108 -1362240 44130 -1362040
rect 44136 -1362240 44158 -1362040
rect 44309 -1362240 44336 -1362040
rect 44337 -1362240 44364 -1362040
rect 44515 -1362240 44537 -1362040
rect 44543 -1362240 44565 -1362040
rect 44716 -1362240 44743 -1362040
rect 44744 -1362240 44771 -1362040
rect 44922 -1362240 44944 -1362040
rect 44950 -1362240 44972 -1362040
rect 45123 -1362240 45150 -1362040
rect 45151 -1362240 45178 -1362040
rect 45329 -1362240 45351 -1362040
rect 45357 -1362240 45379 -1362040
rect 45530 -1362240 45557 -1362040
rect 45558 -1362240 45585 -1362040
rect 45736 -1362240 45758 -1362040
rect 45764 -1362240 45786 -1362040
rect 45937 -1362240 45964 -1362040
rect 45965 -1362240 45992 -1362040
rect 46143 -1362240 46165 -1362040
rect 46171 -1362240 46193 -1362040
rect 46344 -1362240 46371 -1362040
rect 46372 -1362240 46399 -1362040
rect 46550 -1362240 46572 -1362040
rect 46578 -1362240 46600 -1362040
rect 46751 -1362240 46778 -1362040
rect 46779 -1362240 46806 -1362040
rect 46957 -1362240 46979 -1362040
rect 46985 -1362240 47007 -1362040
rect 47158 -1362240 47185 -1362040
rect 47186 -1362240 47213 -1362040
rect 47364 -1362240 47386 -1362040
rect 47392 -1362240 47414 -1362040
rect 47565 -1362240 47592 -1362040
rect 47593 -1362240 47620 -1362040
rect 47771 -1362240 47793 -1362040
rect 47799 -1362240 47821 -1362040
rect 47972 -1362240 47999 -1362040
rect 48000 -1362240 48027 -1362040
rect 48178 -1362240 48200 -1362040
rect 48206 -1362240 48228 -1362040
rect 48379 -1362240 48406 -1362040
rect 48407 -1362240 48434 -1362040
rect 48585 -1362240 48607 -1362040
rect 48613 -1362240 48635 -1362040
rect 48786 -1362240 48813 -1362040
rect 48814 -1362240 48841 -1362040
rect 48992 -1362240 49014 -1362040
rect 49020 -1362240 49042 -1362040
rect 49193 -1362240 49220 -1362040
rect 49221 -1362240 49248 -1362040
rect 49399 -1362240 49421 -1362040
rect 49427 -1362240 49449 -1362040
rect 49600 -1362240 49627 -1362040
rect 49628 -1362240 49655 -1362040
rect 49806 -1362240 49828 -1362040
rect 49834 -1362240 49856 -1362040
rect 50007 -1362240 50034 -1362040
rect 50035 -1362240 50062 -1362040
rect 50213 -1362240 50235 -1362040
rect 50241 -1362240 50263 -1362040
rect 50414 -1362240 50441 -1362040
rect 50442 -1362240 50469 -1362040
rect 50620 -1362240 50642 -1362040
rect 50648 -1362240 50670 -1362040
rect 50821 -1362240 50848 -1362040
rect 50849 -1362240 50876 -1362040
rect 51027 -1362240 51049 -1362040
rect 51055 -1362240 51077 -1362040
rect 51228 -1362240 51255 -1362040
rect 51256 -1362240 51283 -1362040
rect 51434 -1362240 51456 -1362040
rect 51462 -1362240 51484 -1362040
rect 51635 -1362240 51662 -1362040
rect 51663 -1362240 51690 -1362040
rect 51841 -1362240 51863 -1362040
rect 51869 -1362240 51891 -1362040
rect 52042 -1362240 52069 -1362040
rect 52070 -1362240 52097 -1362040
rect 52248 -1362240 52270 -1362040
rect 52276 -1362240 52298 -1362040
rect 52449 -1362240 52476 -1362040
rect 52477 -1362240 52504 -1362040
rect 52655 -1362240 52677 -1362040
rect 52683 -1362240 52705 -1362040
rect 52856 -1362240 52883 -1362040
rect 52884 -1362240 52911 -1362040
rect 53062 -1362240 53084 -1362040
rect 53090 -1362240 53112 -1362040
rect 53263 -1362240 53290 -1362040
rect 53291 -1362240 53318 -1362040
rect 53469 -1362240 53491 -1362040
rect 53497 -1362240 53519 -1362040
rect 53670 -1362240 53697 -1362040
rect 53698 -1362240 53725 -1362040
rect 53876 -1362240 53898 -1362040
rect 53904 -1362240 53926 -1362040
rect 38410 -1362640 38432 -1362440
rect 38438 -1362640 38460 -1362440
rect 38611 -1362640 38638 -1362440
rect 38639 -1362640 38666 -1362440
rect 38812 -1362640 38839 -1362440
rect 38840 -1362640 38867 -1362440
rect 39013 -1362640 39040 -1362440
rect 39041 -1362640 39068 -1362440
rect 39219 -1362640 39241 -1362440
rect 39247 -1362640 39269 -1362440
rect 39425 -1362640 39447 -1362440
rect 39453 -1362640 39475 -1362440
rect 39626 -1362640 39653 -1362440
rect 39654 -1362640 39681 -1362440
rect 39827 -1362640 39854 -1362440
rect 39855 -1362640 39882 -1362440
rect 40033 -1362640 40055 -1362440
rect 40061 -1362640 40083 -1362440
rect 40239 -1362640 40261 -1362440
rect 40267 -1362640 40289 -1362440
rect 40445 -1362640 40467 -1362440
rect 40473 -1362640 40495 -1362440
rect 40646 -1362640 40673 -1362440
rect 40674 -1362640 40701 -1362440
rect 40852 -1362640 40874 -1362440
rect 40880 -1362640 40902 -1362440
rect 41053 -1362640 41080 -1362440
rect 41081 -1362640 41108 -1362440
rect 41259 -1362640 41281 -1362440
rect 41287 -1362640 41309 -1362440
rect 41460 -1362640 41487 -1362440
rect 41488 -1362640 41515 -1362440
rect 41666 -1362640 41688 -1362440
rect 41694 -1362640 41716 -1362440
rect 41867 -1362640 41894 -1362440
rect 41895 -1362640 41922 -1362440
rect 42073 -1362640 42095 -1362440
rect 42101 -1362640 42123 -1362440
rect 42274 -1362640 42301 -1362440
rect 42302 -1362640 42329 -1362440
rect 42480 -1362640 42502 -1362440
rect 42508 -1362640 42530 -1362440
rect 42686 -1362640 42708 -1362440
rect 42714 -1362640 42736 -1362440
rect 42887 -1362640 42914 -1362440
rect 42915 -1362640 42942 -1362440
rect 43088 -1362640 43115 -1362440
rect 43116 -1362640 43143 -1362440
rect 43294 -1362640 43316 -1362440
rect 43322 -1362640 43344 -1362440
rect 43495 -1362640 43522 -1362440
rect 43523 -1362640 43550 -1362440
rect 43701 -1362640 43723 -1362440
rect 43729 -1362640 43751 -1362440
rect 43902 -1362640 43929 -1362440
rect 43930 -1362640 43957 -1362440
rect 44108 -1362640 44130 -1362440
rect 44136 -1362640 44158 -1362440
rect 44309 -1362640 44336 -1362440
rect 44337 -1362640 44364 -1362440
rect 44515 -1362640 44537 -1362440
rect 44543 -1362640 44565 -1362440
rect 44716 -1362640 44743 -1362440
rect 44744 -1362640 44771 -1362440
rect 44922 -1362640 44944 -1362440
rect 44950 -1362640 44972 -1362440
rect 45123 -1362640 45150 -1362440
rect 45151 -1362640 45178 -1362440
rect 45329 -1362640 45351 -1362440
rect 45357 -1362640 45379 -1362440
rect 45530 -1362640 45557 -1362440
rect 45558 -1362640 45585 -1362440
rect 45736 -1362640 45758 -1362440
rect 45764 -1362640 45786 -1362440
rect 45937 -1362640 45964 -1362440
rect 45965 -1362640 45992 -1362440
rect 46143 -1362640 46165 -1362440
rect 46171 -1362640 46193 -1362440
rect 46344 -1362640 46371 -1362440
rect 46372 -1362640 46399 -1362440
rect 46550 -1362640 46572 -1362440
rect 46578 -1362640 46600 -1362440
rect 46751 -1362640 46778 -1362440
rect 46779 -1362640 46806 -1362440
rect 46957 -1362640 46979 -1362440
rect 46985 -1362640 47007 -1362440
rect 47158 -1362640 47185 -1362440
rect 47186 -1362640 47213 -1362440
rect 47364 -1362640 47386 -1362440
rect 47392 -1362640 47414 -1362440
rect 47565 -1362640 47592 -1362440
rect 47593 -1362640 47620 -1362440
rect 47771 -1362640 47793 -1362440
rect 47799 -1362640 47821 -1362440
rect 47972 -1362640 47999 -1362440
rect 48000 -1362640 48027 -1362440
rect 48178 -1362640 48200 -1362440
rect 48206 -1362640 48228 -1362440
rect 48379 -1362640 48406 -1362440
rect 48407 -1362640 48434 -1362440
rect 48585 -1362640 48607 -1362440
rect 48613 -1362640 48635 -1362440
rect 48786 -1362640 48813 -1362440
rect 48814 -1362640 48841 -1362440
rect 48992 -1362640 49014 -1362440
rect 49020 -1362640 49042 -1362440
rect 49193 -1362640 49220 -1362440
rect 49221 -1362640 49248 -1362440
rect 49399 -1362640 49421 -1362440
rect 49427 -1362640 49449 -1362440
rect 49600 -1362640 49627 -1362440
rect 49628 -1362640 49655 -1362440
rect 49806 -1362640 49828 -1362440
rect 49834 -1362640 49856 -1362440
rect 50007 -1362640 50034 -1362440
rect 50035 -1362640 50062 -1362440
rect 50213 -1362640 50235 -1362440
rect 50241 -1362640 50263 -1362440
rect 50414 -1362640 50441 -1362440
rect 50442 -1362640 50469 -1362440
rect 50620 -1362640 50642 -1362440
rect 50648 -1362640 50670 -1362440
rect 50821 -1362640 50848 -1362440
rect 50849 -1362640 50876 -1362440
rect 51027 -1362640 51049 -1362440
rect 51055 -1362640 51077 -1362440
rect 51228 -1362640 51255 -1362440
rect 51256 -1362640 51283 -1362440
rect 51434 -1362640 51456 -1362440
rect 51462 -1362640 51484 -1362440
rect 51635 -1362640 51662 -1362440
rect 51663 -1362640 51690 -1362440
rect 51841 -1362640 51863 -1362440
rect 51869 -1362640 51891 -1362440
rect 52042 -1362640 52069 -1362440
rect 52070 -1362640 52097 -1362440
rect 52248 -1362640 52270 -1362440
rect 52276 -1362640 52298 -1362440
rect 52449 -1362640 52476 -1362440
rect 52477 -1362640 52504 -1362440
rect 52655 -1362640 52677 -1362440
rect 52683 -1362640 52705 -1362440
rect 52856 -1362640 52883 -1362440
rect 52884 -1362640 52911 -1362440
rect 53062 -1362640 53084 -1362440
rect 53090 -1362640 53112 -1362440
rect 53263 -1362640 53290 -1362440
rect 53291 -1362640 53318 -1362440
rect 53469 -1362640 53491 -1362440
rect 53497 -1362640 53519 -1362440
rect 53670 -1362640 53697 -1362440
rect 53698 -1362640 53725 -1362440
rect 53876 -1362640 53898 -1362440
rect 53904 -1362640 53926 -1362440
rect 38611 -1363040 38638 -1362840
rect 38639 -1363040 38666 -1362840
rect 38812 -1363040 38839 -1362840
rect 38840 -1363040 38867 -1362840
rect 39013 -1363040 39040 -1362840
rect 39041 -1363040 39068 -1362840
rect 39219 -1363040 39241 -1362840
rect 39247 -1363040 39269 -1362840
rect 39425 -1363040 39447 -1362840
rect 39453 -1363040 39475 -1362840
rect 39626 -1363040 39653 -1362840
rect 39654 -1363040 39681 -1362840
rect 39827 -1363040 39854 -1362840
rect 39855 -1363040 39882 -1362840
rect 40033 -1363040 40055 -1362840
rect 40061 -1363040 40083 -1362840
rect 40239 -1363040 40261 -1362840
rect 40267 -1363040 40289 -1362840
rect 40445 -1363040 40467 -1362840
rect 40473 -1363040 40495 -1362840
rect 40646 -1363040 40673 -1362840
rect 40674 -1363040 40701 -1362840
rect 40852 -1363040 40874 -1362840
rect 40880 -1363040 40902 -1362840
rect 41053 -1363040 41080 -1362840
rect 41081 -1363040 41108 -1362840
rect 41259 -1363040 41281 -1362840
rect 41287 -1363040 41309 -1362840
rect 41460 -1363040 41487 -1362840
rect 41488 -1363040 41515 -1362840
rect 41666 -1363040 41688 -1362840
rect 41694 -1363040 41716 -1362840
rect 41867 -1363040 41894 -1362840
rect 41895 -1363040 41922 -1362840
rect 42073 -1363040 42095 -1362840
rect 42101 -1363040 42123 -1362840
rect 42274 -1363040 42301 -1362840
rect 42302 -1363040 42329 -1362840
rect 42480 -1363040 42502 -1362840
rect 42508 -1363040 42530 -1362840
rect 42686 -1363040 42708 -1362840
rect 42714 -1363040 42736 -1362840
rect 42887 -1363040 42914 -1362840
rect 42915 -1363040 42942 -1362840
rect 43088 -1363040 43115 -1362840
rect 43116 -1363040 43143 -1362840
rect 43294 -1363040 43316 -1362840
rect 43322 -1363040 43344 -1362840
rect 43495 -1363040 43522 -1362840
rect 43523 -1363040 43550 -1362840
rect 43701 -1363040 43723 -1362840
rect 43729 -1363040 43751 -1362840
rect 43902 -1363040 43929 -1362840
rect 43930 -1363040 43957 -1362840
rect 44108 -1363040 44130 -1362840
rect 44136 -1363040 44158 -1362840
rect 44309 -1363040 44336 -1362840
rect 44337 -1363040 44364 -1362840
rect 44515 -1363040 44537 -1362840
rect 44543 -1363040 44565 -1362840
rect 44716 -1363040 44743 -1362840
rect 44744 -1363040 44771 -1362840
rect 44922 -1363040 44944 -1362840
rect 44950 -1363040 44972 -1362840
rect 45123 -1363040 45150 -1362840
rect 45151 -1363040 45178 -1362840
rect 45329 -1363040 45351 -1362840
rect 45357 -1363040 45379 -1362840
rect 45530 -1363040 45557 -1362840
rect 45558 -1363040 45585 -1362840
rect 45736 -1363040 45758 -1362840
rect 45764 -1363040 45786 -1362840
rect 45937 -1363040 45964 -1362840
rect 45965 -1363040 45992 -1362840
rect 46143 -1363040 46165 -1362840
rect 46171 -1363040 46193 -1362840
rect 46344 -1363040 46371 -1362840
rect 46372 -1363040 46399 -1362840
rect 46550 -1363040 46572 -1362840
rect 46578 -1363040 46600 -1362840
rect 46751 -1363040 46778 -1362840
rect 46779 -1363040 46806 -1362840
rect 46957 -1363040 46979 -1362840
rect 46985 -1363040 47007 -1362840
rect 47158 -1363040 47185 -1362840
rect 47186 -1363040 47213 -1362840
rect 47364 -1363040 47386 -1362840
rect 47392 -1363040 47414 -1362840
rect 47565 -1363040 47592 -1362840
rect 47593 -1363040 47620 -1362840
rect 47771 -1363040 47793 -1362840
rect 47799 -1363040 47821 -1362840
rect 47972 -1363040 47999 -1362840
rect 48000 -1363040 48027 -1362840
rect 48178 -1363040 48200 -1362840
rect 48206 -1363040 48228 -1362840
rect 48379 -1363040 48406 -1362840
rect 48407 -1363040 48434 -1362840
rect 48585 -1363040 48607 -1362840
rect 48613 -1363040 48635 -1362840
rect 48786 -1363040 48813 -1362840
rect 48814 -1363040 48841 -1362840
rect 48992 -1363040 49014 -1362840
rect 49020 -1363040 49042 -1362840
rect 49193 -1363040 49220 -1362840
rect 49221 -1363040 49248 -1362840
rect 49399 -1363040 49421 -1362840
rect 49427 -1363040 49449 -1362840
rect 49600 -1363040 49627 -1362840
rect 49628 -1363040 49655 -1362840
rect 49806 -1363040 49828 -1362840
rect 49834 -1363040 49856 -1362840
rect 50007 -1363040 50034 -1362840
rect 50035 -1363040 50062 -1362840
rect 50213 -1363040 50235 -1362840
rect 50241 -1363040 50263 -1362840
rect 50414 -1363040 50441 -1362840
rect 50442 -1363040 50469 -1362840
rect 50620 -1363040 50642 -1362840
rect 50648 -1363040 50670 -1362840
rect 50821 -1363040 50848 -1362840
rect 50849 -1363040 50876 -1362840
rect 51027 -1363040 51049 -1362840
rect 51055 -1363040 51077 -1362840
rect 51228 -1363040 51255 -1362840
rect 51256 -1363040 51283 -1362840
rect 51434 -1363040 51456 -1362840
rect 51462 -1363040 51484 -1362840
rect 51635 -1363040 51662 -1362840
rect 51663 -1363040 51690 -1362840
rect 51841 -1363040 51863 -1362840
rect 51869 -1363040 51891 -1362840
rect 52042 -1363040 52069 -1362840
rect 52070 -1363040 52097 -1362840
rect 52248 -1363040 52270 -1362840
rect 52276 -1363040 52298 -1362840
rect 52449 -1363040 52476 -1362840
rect 52477 -1363040 52504 -1362840
rect 52655 -1363040 52677 -1362840
rect 52683 -1363040 52705 -1362840
rect 52856 -1363040 52883 -1362840
rect 52884 -1363040 52911 -1362840
rect 53062 -1363040 53084 -1362840
rect 53090 -1363040 53112 -1362840
rect 53263 -1363040 53290 -1362840
rect 53291 -1363040 53318 -1362840
rect 53469 -1363040 53491 -1362840
rect 53497 -1363040 53519 -1362840
rect 53670 -1363040 53697 -1362840
rect 53698 -1363040 53725 -1362840
rect 53876 -1363040 53898 -1362840
rect 53904 -1363040 53926 -1362840
rect 38611 -1363440 38638 -1363240
rect 38639 -1363440 38666 -1363240
rect 38812 -1363440 38839 -1363240
rect 38840 -1363440 38867 -1363240
rect 39013 -1363440 39040 -1363240
rect 39041 -1363440 39068 -1363240
rect 39219 -1363440 39241 -1363240
rect 39247 -1363440 39269 -1363240
rect 39425 -1363440 39447 -1363240
rect 39453 -1363440 39475 -1363240
rect 39626 -1363440 39653 -1363240
rect 39654 -1363440 39681 -1363240
rect 39827 -1363440 39854 -1363240
rect 39855 -1363440 39882 -1363240
rect 40033 -1363440 40055 -1363240
rect 40061 -1363440 40083 -1363240
rect 40239 -1363440 40261 -1363240
rect 40267 -1363440 40289 -1363240
rect 40445 -1363440 40467 -1363240
rect 40473 -1363440 40495 -1363240
rect 40646 -1363440 40673 -1363240
rect 40674 -1363440 40701 -1363240
rect 40852 -1363440 40874 -1363240
rect 40880 -1363440 40902 -1363240
rect 41053 -1363440 41080 -1363240
rect 41081 -1363440 41108 -1363240
rect 41259 -1363440 41281 -1363240
rect 41287 -1363440 41309 -1363240
rect 41460 -1363440 41487 -1363240
rect 41488 -1363440 41515 -1363240
rect 41666 -1363440 41688 -1363240
rect 41694 -1363440 41716 -1363240
rect 41867 -1363440 41894 -1363240
rect 41895 -1363440 41922 -1363240
rect 42073 -1363440 42095 -1363240
rect 42101 -1363440 42123 -1363240
rect 42274 -1363440 42301 -1363240
rect 42302 -1363440 42329 -1363240
rect 42480 -1363440 42502 -1363240
rect 42508 -1363440 42530 -1363240
rect 42686 -1363440 42708 -1363240
rect 42714 -1363440 42736 -1363240
rect 42887 -1363440 42914 -1363240
rect 42915 -1363440 42942 -1363240
rect 43088 -1363440 43115 -1363240
rect 43116 -1363440 43143 -1363240
rect 43294 -1363440 43316 -1363240
rect 43322 -1363440 43344 -1363240
rect 43495 -1363440 43522 -1363240
rect 43523 -1363440 43550 -1363240
rect 43701 -1363440 43723 -1363240
rect 43729 -1363440 43751 -1363240
rect 43902 -1363440 43929 -1363240
rect 43930 -1363440 43957 -1363240
rect 44108 -1363440 44130 -1363240
rect 44136 -1363440 44158 -1363240
rect 44309 -1363440 44336 -1363240
rect 44337 -1363440 44364 -1363240
rect 44515 -1363440 44537 -1363240
rect 44543 -1363440 44565 -1363240
rect 44716 -1363440 44743 -1363240
rect 44744 -1363440 44771 -1363240
rect 44922 -1363440 44944 -1363240
rect 44950 -1363440 44972 -1363240
rect 45123 -1363440 45150 -1363240
rect 45151 -1363440 45178 -1363240
rect 45329 -1363440 45351 -1363240
rect 45357 -1363440 45379 -1363240
rect 45530 -1363440 45557 -1363240
rect 45558 -1363440 45585 -1363240
rect 45736 -1363440 45758 -1363240
rect 45764 -1363440 45786 -1363240
rect 45937 -1363440 45964 -1363240
rect 45965 -1363440 45992 -1363240
rect 46143 -1363440 46165 -1363240
rect 46171 -1363440 46193 -1363240
rect 46344 -1363440 46371 -1363240
rect 46372 -1363440 46399 -1363240
rect 46550 -1363440 46572 -1363240
rect 46578 -1363440 46600 -1363240
rect 46751 -1363440 46778 -1363240
rect 46779 -1363440 46806 -1363240
rect 46957 -1363440 46979 -1363240
rect 46985 -1363440 47007 -1363240
rect 47158 -1363440 47185 -1363240
rect 47186 -1363440 47213 -1363240
rect 47364 -1363440 47386 -1363240
rect 47392 -1363440 47414 -1363240
rect 47565 -1363440 47592 -1363240
rect 47593 -1363440 47620 -1363240
rect 47771 -1363440 47793 -1363240
rect 47799 -1363440 47821 -1363240
rect 47972 -1363440 47999 -1363240
rect 48000 -1363440 48027 -1363240
rect 48178 -1363440 48200 -1363240
rect 48206 -1363440 48228 -1363240
rect 48379 -1363440 48406 -1363240
rect 48407 -1363440 48434 -1363240
rect 48585 -1363440 48607 -1363240
rect 48613 -1363440 48635 -1363240
rect 48786 -1363440 48813 -1363240
rect 48814 -1363440 48841 -1363240
rect 48992 -1363440 49014 -1363240
rect 49020 -1363440 49042 -1363240
rect 49193 -1363440 49220 -1363240
rect 49221 -1363440 49248 -1363240
rect 49399 -1363440 49421 -1363240
rect 49427 -1363440 49449 -1363240
rect 49600 -1363440 49627 -1363240
rect 49628 -1363440 49655 -1363240
rect 49806 -1363440 49828 -1363240
rect 49834 -1363440 49856 -1363240
rect 50007 -1363440 50034 -1363240
rect 50035 -1363440 50062 -1363240
rect 50213 -1363440 50235 -1363240
rect 50241 -1363440 50263 -1363240
rect 50414 -1363440 50441 -1363240
rect 50442 -1363440 50469 -1363240
rect 50620 -1363440 50642 -1363240
rect 50648 -1363440 50670 -1363240
rect 50821 -1363440 50848 -1363240
rect 50849 -1363440 50876 -1363240
rect 51027 -1363440 51049 -1363240
rect 51055 -1363440 51077 -1363240
rect 51228 -1363440 51255 -1363240
rect 51256 -1363440 51283 -1363240
rect 51434 -1363440 51456 -1363240
rect 51462 -1363440 51484 -1363240
rect 51635 -1363440 51662 -1363240
rect 51663 -1363440 51690 -1363240
rect 51841 -1363440 51863 -1363240
rect 51869 -1363440 51891 -1363240
rect 52042 -1363440 52069 -1363240
rect 52070 -1363440 52097 -1363240
rect 52248 -1363440 52270 -1363240
rect 52276 -1363440 52298 -1363240
rect 52449 -1363440 52476 -1363240
rect 52477 -1363440 52504 -1363240
rect 52655 -1363440 52677 -1363240
rect 52683 -1363440 52705 -1363240
rect 52856 -1363440 52883 -1363240
rect 52884 -1363440 52911 -1363240
rect 53062 -1363440 53084 -1363240
rect 53090 -1363440 53112 -1363240
rect 53263 -1363440 53290 -1363240
rect 53291 -1363440 53318 -1363240
rect 53469 -1363440 53491 -1363240
rect 53497 -1363440 53519 -1363240
rect 53670 -1363440 53697 -1363240
rect 53698 -1363440 53725 -1363240
rect 53876 -1363440 53898 -1363240
rect 53904 -1363440 53926 -1363240
rect 38611 -1363840 38638 -1363640
rect 38639 -1363840 38666 -1363640
rect 38812 -1363840 38839 -1363640
rect 38840 -1363840 38867 -1363640
rect 39013 -1363840 39040 -1363640
rect 39041 -1363840 39068 -1363640
rect 39219 -1363840 39241 -1363640
rect 39247 -1363840 39269 -1363640
rect 39425 -1363840 39447 -1363640
rect 39453 -1363840 39475 -1363640
rect 39626 -1363840 39653 -1363640
rect 39654 -1363840 39681 -1363640
rect 39827 -1363840 39854 -1363640
rect 39855 -1363840 39882 -1363640
rect 40033 -1363840 40055 -1363640
rect 40061 -1363840 40083 -1363640
rect 40239 -1363840 40261 -1363640
rect 40267 -1363840 40289 -1363640
rect 40445 -1363840 40467 -1363640
rect 40473 -1363840 40495 -1363640
rect 40646 -1363840 40673 -1363640
rect 40674 -1363840 40701 -1363640
rect 40852 -1363840 40874 -1363640
rect 40880 -1363840 40902 -1363640
rect 41053 -1363840 41080 -1363640
rect 41081 -1363840 41108 -1363640
rect 41259 -1363840 41281 -1363640
rect 41287 -1363840 41309 -1363640
rect 41460 -1363840 41487 -1363640
rect 41488 -1363840 41515 -1363640
rect 41666 -1363840 41688 -1363640
rect 41694 -1363840 41716 -1363640
rect 41867 -1363840 41894 -1363640
rect 41895 -1363840 41922 -1363640
rect 42073 -1363840 42095 -1363640
rect 42101 -1363840 42123 -1363640
rect 42274 -1363840 42301 -1363640
rect 42302 -1363840 42329 -1363640
rect 42480 -1363840 42502 -1363640
rect 42508 -1363840 42530 -1363640
rect 42686 -1363840 42708 -1363640
rect 42714 -1363840 42736 -1363640
rect 42887 -1363840 42914 -1363640
rect 42915 -1363840 42942 -1363640
rect 43088 -1363840 43115 -1363640
rect 43116 -1363840 43143 -1363640
rect 43294 -1363840 43316 -1363640
rect 43322 -1363840 43344 -1363640
rect 43495 -1363840 43522 -1363640
rect 43523 -1363840 43550 -1363640
rect 43701 -1363840 43723 -1363640
rect 43729 -1363840 43751 -1363640
rect 43902 -1363840 43929 -1363640
rect 43930 -1363840 43957 -1363640
rect 44108 -1363840 44130 -1363640
rect 44136 -1363840 44158 -1363640
rect 44309 -1363840 44336 -1363640
rect 44337 -1363840 44364 -1363640
rect 44515 -1363840 44537 -1363640
rect 44543 -1363840 44565 -1363640
rect 44716 -1363840 44743 -1363640
rect 44744 -1363840 44771 -1363640
rect 44922 -1363840 44944 -1363640
rect 44950 -1363840 44972 -1363640
rect 45123 -1363840 45150 -1363640
rect 45151 -1363840 45178 -1363640
rect 45329 -1363840 45351 -1363640
rect 45357 -1363840 45379 -1363640
rect 45530 -1363840 45557 -1363640
rect 45558 -1363840 45585 -1363640
rect 45736 -1363840 45758 -1363640
rect 45764 -1363840 45786 -1363640
rect 45937 -1363840 45964 -1363640
rect 45965 -1363840 45992 -1363640
rect 46143 -1363840 46165 -1363640
rect 46171 -1363840 46193 -1363640
rect 46344 -1363840 46371 -1363640
rect 46372 -1363840 46399 -1363640
rect 46550 -1363840 46572 -1363640
rect 46578 -1363840 46600 -1363640
rect 46751 -1363840 46778 -1363640
rect 46779 -1363840 46806 -1363640
rect 46957 -1363840 46979 -1363640
rect 46985 -1363840 47007 -1363640
rect 47158 -1363840 47185 -1363640
rect 47186 -1363840 47213 -1363640
rect 47364 -1363840 47386 -1363640
rect 47392 -1363840 47414 -1363640
rect 47565 -1363840 47592 -1363640
rect 47593 -1363840 47620 -1363640
rect 47771 -1363840 47793 -1363640
rect 47799 -1363840 47821 -1363640
rect 47972 -1363840 47999 -1363640
rect 48000 -1363840 48027 -1363640
rect 48178 -1363840 48200 -1363640
rect 48206 -1363840 48228 -1363640
rect 48379 -1363840 48406 -1363640
rect 48407 -1363840 48434 -1363640
rect 48585 -1363840 48607 -1363640
rect 48613 -1363840 48635 -1363640
rect 48786 -1363840 48813 -1363640
rect 48814 -1363840 48841 -1363640
rect 48992 -1363840 49014 -1363640
rect 49020 -1363840 49042 -1363640
rect 49193 -1363840 49220 -1363640
rect 49221 -1363840 49248 -1363640
rect 49399 -1363840 49421 -1363640
rect 49427 -1363840 49449 -1363640
rect 49600 -1363840 49627 -1363640
rect 49628 -1363840 49655 -1363640
rect 49806 -1363840 49828 -1363640
rect 49834 -1363840 49856 -1363640
rect 50007 -1363840 50034 -1363640
rect 50035 -1363840 50062 -1363640
rect 50213 -1363840 50235 -1363640
rect 50241 -1363840 50263 -1363640
rect 50414 -1363840 50441 -1363640
rect 50442 -1363840 50469 -1363640
rect 50620 -1363840 50642 -1363640
rect 50648 -1363840 50670 -1363640
rect 50821 -1363840 50848 -1363640
rect 50849 -1363840 50876 -1363640
rect 51027 -1363840 51049 -1363640
rect 51055 -1363840 51077 -1363640
rect 51228 -1363840 51255 -1363640
rect 51256 -1363840 51283 -1363640
rect 51434 -1363840 51456 -1363640
rect 51462 -1363840 51484 -1363640
rect 51635 -1363840 51662 -1363640
rect 51663 -1363840 51690 -1363640
rect 51841 -1363840 51863 -1363640
rect 51869 -1363840 51891 -1363640
rect 52042 -1363840 52069 -1363640
rect 52070 -1363840 52097 -1363640
rect 52248 -1363840 52270 -1363640
rect 52276 -1363840 52298 -1363640
rect 52449 -1363840 52476 -1363640
rect 52477 -1363840 52504 -1363640
rect 52655 -1363840 52677 -1363640
rect 52683 -1363840 52705 -1363640
rect 52856 -1363840 52883 -1363640
rect 52884 -1363840 52911 -1363640
rect 53062 -1363840 53084 -1363640
rect 53090 -1363840 53112 -1363640
rect 53263 -1363840 53290 -1363640
rect 53291 -1363840 53318 -1363640
rect 53469 -1363840 53491 -1363640
rect 53497 -1363840 53519 -1363640
rect 53670 -1363840 53697 -1363640
rect 53698 -1363840 53725 -1363640
rect 53876 -1363840 53898 -1363640
rect 53904 -1363840 53926 -1363640
rect 38611 -1364240 38638 -1364040
rect 38639 -1364240 38666 -1364040
rect 38812 -1364240 38839 -1364040
rect 38840 -1364240 38867 -1364040
rect 39013 -1364240 39040 -1364040
rect 39041 -1364240 39068 -1364040
rect 39219 -1364240 39241 -1364040
rect 39247 -1364240 39269 -1364040
rect 39425 -1364240 39447 -1364040
rect 39453 -1364240 39475 -1364040
rect 39626 -1364240 39653 -1364040
rect 39654 -1364240 39681 -1364040
rect 39827 -1364240 39854 -1364040
rect 39855 -1364240 39882 -1364040
rect 40033 -1364240 40055 -1364040
rect 40061 -1364240 40083 -1364040
rect 40239 -1364240 40261 -1364040
rect 40267 -1364240 40289 -1364040
rect 40445 -1364240 40467 -1364040
rect 40473 -1364240 40495 -1364040
rect 40646 -1364240 40673 -1364040
rect 40674 -1364240 40701 -1364040
rect 40852 -1364240 40874 -1364040
rect 40880 -1364240 40902 -1364040
rect 41053 -1364240 41080 -1364040
rect 41081 -1364240 41108 -1364040
rect 41259 -1364240 41281 -1364040
rect 41287 -1364240 41309 -1364040
rect 41460 -1364240 41487 -1364040
rect 41488 -1364240 41515 -1364040
rect 41666 -1364240 41688 -1364040
rect 41694 -1364240 41716 -1364040
rect 41867 -1364240 41894 -1364040
rect 41895 -1364240 41922 -1364040
rect 42073 -1364240 42095 -1364040
rect 42101 -1364240 42123 -1364040
rect 42274 -1364240 42301 -1364040
rect 42302 -1364240 42329 -1364040
rect 42480 -1364240 42502 -1364040
rect 42508 -1364240 42530 -1364040
rect 42686 -1364240 42708 -1364040
rect 42714 -1364240 42736 -1364040
rect 42887 -1364240 42914 -1364040
rect 42915 -1364240 42942 -1364040
rect 43088 -1364240 43115 -1364040
rect 43116 -1364240 43143 -1364040
rect 43294 -1364240 43316 -1364040
rect 43322 -1364240 43344 -1364040
rect 43495 -1364240 43522 -1364040
rect 43523 -1364240 43550 -1364040
rect 43701 -1364240 43723 -1364040
rect 43729 -1364240 43751 -1364040
rect 43902 -1364240 43929 -1364040
rect 43930 -1364240 43957 -1364040
rect 44108 -1364240 44130 -1364040
rect 44136 -1364240 44158 -1364040
rect 44309 -1364240 44336 -1364040
rect 44337 -1364240 44364 -1364040
rect 44515 -1364240 44537 -1364040
rect 44543 -1364240 44565 -1364040
rect 44716 -1364240 44743 -1364040
rect 44744 -1364240 44771 -1364040
rect 44922 -1364240 44944 -1364040
rect 44950 -1364240 44972 -1364040
rect 45123 -1364240 45150 -1364040
rect 45151 -1364240 45178 -1364040
rect 45329 -1364240 45351 -1364040
rect 45357 -1364240 45379 -1364040
rect 45530 -1364240 45557 -1364040
rect 45558 -1364240 45585 -1364040
rect 45736 -1364240 45758 -1364040
rect 45764 -1364240 45786 -1364040
rect 45937 -1364240 45964 -1364040
rect 45965 -1364240 45992 -1364040
rect 46143 -1364240 46165 -1364040
rect 46171 -1364240 46193 -1364040
rect 46344 -1364240 46371 -1364040
rect 46372 -1364240 46399 -1364040
rect 46550 -1364240 46572 -1364040
rect 46578 -1364240 46600 -1364040
rect 46751 -1364240 46778 -1364040
rect 46779 -1364240 46806 -1364040
rect 46957 -1364240 46979 -1364040
rect 46985 -1364240 47007 -1364040
rect 47158 -1364240 47185 -1364040
rect 47186 -1364240 47213 -1364040
rect 47364 -1364240 47386 -1364040
rect 47392 -1364240 47414 -1364040
rect 47565 -1364240 47592 -1364040
rect 47593 -1364240 47620 -1364040
rect 47771 -1364240 47793 -1364040
rect 47799 -1364240 47821 -1364040
rect 47972 -1364240 47999 -1364040
rect 48000 -1364240 48027 -1364040
rect 48178 -1364240 48200 -1364040
rect 48206 -1364240 48228 -1364040
rect 48379 -1364240 48406 -1364040
rect 48407 -1364240 48434 -1364040
rect 48585 -1364240 48607 -1364040
rect 48613 -1364240 48635 -1364040
rect 48786 -1364240 48813 -1364040
rect 48814 -1364240 48841 -1364040
rect 48992 -1364240 49014 -1364040
rect 49020 -1364240 49042 -1364040
rect 49193 -1364240 49220 -1364040
rect 49221 -1364240 49248 -1364040
rect 49399 -1364240 49421 -1364040
rect 49427 -1364240 49449 -1364040
rect 49600 -1364240 49627 -1364040
rect 49628 -1364240 49655 -1364040
rect 49806 -1364240 49828 -1364040
rect 49834 -1364240 49856 -1364040
rect 50007 -1364240 50034 -1364040
rect 50035 -1364240 50062 -1364040
rect 50213 -1364240 50235 -1364040
rect 50241 -1364240 50263 -1364040
rect 50414 -1364240 50441 -1364040
rect 50442 -1364240 50469 -1364040
rect 50620 -1364240 50642 -1364040
rect 50648 -1364240 50670 -1364040
rect 50821 -1364240 50848 -1364040
rect 50849 -1364240 50876 -1364040
rect 51027 -1364240 51049 -1364040
rect 51055 -1364240 51077 -1364040
rect 51228 -1364240 51255 -1364040
rect 51256 -1364240 51283 -1364040
rect 51434 -1364240 51456 -1364040
rect 51462 -1364240 51484 -1364040
rect 51635 -1364240 51662 -1364040
rect 51663 -1364240 51690 -1364040
rect 51841 -1364240 51863 -1364040
rect 51869 -1364240 51891 -1364040
rect 52042 -1364240 52069 -1364040
rect 52070 -1364240 52097 -1364040
rect 52248 -1364240 52270 -1364040
rect 52276 -1364240 52298 -1364040
rect 52449 -1364240 52476 -1364040
rect 52477 -1364240 52504 -1364040
rect 52655 -1364240 52677 -1364040
rect 52683 -1364240 52705 -1364040
rect 52856 -1364240 52883 -1364040
rect 52884 -1364240 52911 -1364040
rect 53062 -1364240 53084 -1364040
rect 53090 -1364240 53112 -1364040
rect 53263 -1364240 53290 -1364040
rect 53291 -1364240 53318 -1364040
rect 53469 -1364240 53491 -1364040
rect 53497 -1364240 53519 -1364040
rect 53670 -1364240 53697 -1364040
rect 53698 -1364240 53725 -1364040
rect 53876 -1364240 53898 -1364040
rect 53904 -1364240 53926 -1364040
rect 38611 -1364640 38638 -1364440
rect 38639 -1364640 38666 -1364440
rect 38812 -1364640 38839 -1364440
rect 38840 -1364640 38867 -1364440
rect 39013 -1364640 39040 -1364440
rect 39041 -1364640 39068 -1364440
rect 39219 -1364640 39241 -1364440
rect 39247 -1364640 39269 -1364440
rect 39425 -1364640 39447 -1364440
rect 39453 -1364640 39475 -1364440
rect 39626 -1364640 39653 -1364440
rect 39654 -1364640 39681 -1364440
rect 39827 -1364640 39854 -1364440
rect 39855 -1364640 39882 -1364440
rect 40033 -1364640 40055 -1364440
rect 40061 -1364640 40083 -1364440
rect 40239 -1364640 40261 -1364440
rect 40267 -1364640 40289 -1364440
rect 40445 -1364640 40467 -1364440
rect 40473 -1364640 40495 -1364440
rect 40646 -1364640 40673 -1364440
rect 40674 -1364640 40701 -1364440
rect 40852 -1364640 40874 -1364440
rect 40880 -1364640 40902 -1364440
rect 41053 -1364640 41080 -1364440
rect 41081 -1364640 41108 -1364440
rect 41259 -1364640 41281 -1364440
rect 41287 -1364640 41309 -1364440
rect 41460 -1364640 41487 -1364440
rect 41488 -1364640 41515 -1364440
rect 41666 -1364640 41688 -1364440
rect 41694 -1364640 41716 -1364440
rect 41867 -1364640 41894 -1364440
rect 41895 -1364640 41922 -1364440
rect 42073 -1364640 42095 -1364440
rect 42101 -1364640 42123 -1364440
rect 42274 -1364640 42301 -1364440
rect 42302 -1364640 42329 -1364440
rect 42480 -1364640 42502 -1364440
rect 42508 -1364640 42530 -1364440
rect 42686 -1364640 42708 -1364440
rect 42714 -1364640 42736 -1364440
rect 42887 -1364640 42914 -1364440
rect 42915 -1364640 42942 -1364440
rect 43088 -1364640 43115 -1364440
rect 43116 -1364640 43143 -1364440
rect 43294 -1364640 43316 -1364440
rect 43322 -1364640 43344 -1364440
rect 43495 -1364640 43522 -1364440
rect 43523 -1364640 43550 -1364440
rect 43701 -1364640 43723 -1364440
rect 43729 -1364640 43751 -1364440
rect 43902 -1364640 43929 -1364440
rect 43930 -1364640 43957 -1364440
rect 44108 -1364640 44130 -1364440
rect 44136 -1364640 44158 -1364440
rect 44309 -1364640 44336 -1364440
rect 44337 -1364640 44364 -1364440
rect 44515 -1364640 44537 -1364440
rect 44543 -1364640 44565 -1364440
rect 44716 -1364640 44743 -1364440
rect 44744 -1364640 44771 -1364440
rect 44922 -1364640 44944 -1364440
rect 44950 -1364640 44972 -1364440
rect 45123 -1364640 45150 -1364440
rect 45151 -1364640 45178 -1364440
rect 45329 -1364640 45351 -1364440
rect 45357 -1364640 45379 -1364440
rect 45530 -1364640 45557 -1364440
rect 45558 -1364640 45585 -1364440
rect 45736 -1364640 45758 -1364440
rect 45764 -1364640 45786 -1364440
rect 45937 -1364640 45964 -1364440
rect 45965 -1364640 45992 -1364440
rect 46143 -1364640 46165 -1364440
rect 46171 -1364640 46193 -1364440
rect 46344 -1364640 46371 -1364440
rect 46372 -1364640 46399 -1364440
rect 46550 -1364640 46572 -1364440
rect 46578 -1364640 46600 -1364440
rect 46751 -1364640 46778 -1364440
rect 46779 -1364640 46806 -1364440
rect 46957 -1364640 46979 -1364440
rect 46985 -1364640 47007 -1364440
rect 47158 -1364640 47185 -1364440
rect 47186 -1364640 47213 -1364440
rect 47364 -1364640 47386 -1364440
rect 47392 -1364640 47414 -1364440
rect 47565 -1364640 47592 -1364440
rect 47593 -1364640 47620 -1364440
rect 47771 -1364640 47793 -1364440
rect 47799 -1364640 47821 -1364440
rect 47972 -1364640 47999 -1364440
rect 48000 -1364640 48027 -1364440
rect 48178 -1364640 48200 -1364440
rect 48206 -1364640 48228 -1364440
rect 48379 -1364640 48406 -1364440
rect 48407 -1364640 48434 -1364440
rect 48585 -1364640 48607 -1364440
rect 48613 -1364640 48635 -1364440
rect 48786 -1364640 48813 -1364440
rect 48814 -1364640 48841 -1364440
rect 48992 -1364640 49014 -1364440
rect 49020 -1364640 49042 -1364440
rect 49193 -1364640 49220 -1364440
rect 49221 -1364640 49248 -1364440
rect 49399 -1364640 49421 -1364440
rect 49427 -1364640 49449 -1364440
rect 49600 -1364640 49627 -1364440
rect 49628 -1364640 49655 -1364440
rect 49806 -1364640 49828 -1364440
rect 49834 -1364640 49856 -1364440
rect 50007 -1364640 50034 -1364440
rect 50035 -1364640 50062 -1364440
rect 50213 -1364640 50235 -1364440
rect 50241 -1364640 50263 -1364440
rect 50414 -1364640 50441 -1364440
rect 50442 -1364640 50469 -1364440
rect 50620 -1364640 50642 -1364440
rect 50648 -1364640 50670 -1364440
rect 50821 -1364640 50848 -1364440
rect 50849 -1364640 50876 -1364440
rect 51027 -1364640 51049 -1364440
rect 51055 -1364640 51077 -1364440
rect 51228 -1364640 51255 -1364440
rect 51256 -1364640 51283 -1364440
rect 51434 -1364640 51456 -1364440
rect 51462 -1364640 51484 -1364440
rect 51635 -1364640 51662 -1364440
rect 51663 -1364640 51690 -1364440
rect 51841 -1364640 51863 -1364440
rect 51869 -1364640 51891 -1364440
rect 52042 -1364640 52069 -1364440
rect 52070 -1364640 52097 -1364440
rect 52248 -1364640 52270 -1364440
rect 52276 -1364640 52298 -1364440
rect 52449 -1364640 52476 -1364440
rect 52477 -1364640 52504 -1364440
rect 52655 -1364640 52677 -1364440
rect 52683 -1364640 52705 -1364440
rect 52856 -1364640 52883 -1364440
rect 52884 -1364640 52911 -1364440
rect 53062 -1364640 53084 -1364440
rect 53090 -1364640 53112 -1364440
rect 53263 -1364640 53290 -1364440
rect 53291 -1364640 53318 -1364440
rect 53469 -1364640 53491 -1364440
rect 53497 -1364640 53519 -1364440
rect 53670 -1364640 53697 -1364440
rect 53698 -1364640 53725 -1364440
rect 53876 -1364640 53898 -1364440
rect 53904 -1364640 53926 -1364440
rect 468 -1367643 503 -1367609
rect 469 -1367662 503 -1367643
rect 488 -1368057 503 -1367662
rect 522 -1367696 557 -1367662
rect 1007 -1367696 1042 -1367662
rect 522 -1368057 556 -1367696
rect 1008 -1367715 1042 -1367696
rect 522 -1368091 537 -1368057
rect 1027 -1368110 1042 -1367715
rect 1061 -1367749 1096 -1367715
rect 1546 -1367749 1581 -1367715
rect 1061 -1368110 1095 -1367749
rect 1547 -1367768 1581 -1367749
rect 1061 -1368144 1076 -1368110
rect 1566 -1368163 1581 -1367768
rect 1600 -1367802 1635 -1367768
rect 2085 -1367802 2120 -1367768
rect 1600 -1368163 1634 -1367802
rect 2086 -1367821 2120 -1367802
rect 1600 -1368197 1615 -1368163
rect 2105 -1368216 2120 -1367821
rect 2139 -1367855 2174 -1367821
rect 2624 -1367855 2659 -1367821
rect 2139 -1368216 2173 -1367855
rect 2625 -1367874 2659 -1367855
rect 2139 -1368250 2154 -1368216
rect 2644 -1368269 2659 -1367874
rect 2678 -1367908 2713 -1367874
rect 3163 -1367908 3198 -1367874
rect 2678 -1368269 2712 -1367908
rect 3164 -1367927 3198 -1367908
rect 2678 -1368303 2693 -1368269
rect 3183 -1368322 3198 -1367927
rect 3217 -1367961 3252 -1367927
rect 3217 -1368322 3251 -1367961
rect 3217 -1368356 3232 -1368322
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
use CNR_GR06_op_amp  CNR_GR06_op_amp_0
timestamp 1713380705
transform 1 0 38514 0 1 -1362440
box 0 -2800 7251 2767
use CNR_GR06_op_amp  CNR_GR06_op_amp_1
timestamp 1713380705
transform 1 0 0 0 1 -1365240
box 0 -2800 7251 2767
use Non_overlapping_clock  Non_overlapping_clock_0
timestamp 1713380705
transform 1 0 38232 0 1 -1363640
box 0 -1600 16866 4475
use CNR_GR06_op_amp  x2
timestamp 1713380705
transform 1 0 38233 0 1 -1365240
box 0 -2800 7251 2767
use Non_overlapping_clock  x9
timestamp 1713380705
transform 1 0 38232 0 1 -1365240
box 0 -1600 16866 4475
use sky130_fd_pr__cap_mim_m3_1_C8GDQN  XC1
timestamp 0
transform 1 0 3186 0 1 -78520
box -3186 -85320 3186 85320
use sky130_fd_pr__cap_mim_m3_1_CWHDQN  XC2
timestamp 0
transform 1 0 9558 0 1 -290360
box -3186 -132720 3186 132720
use sky130_fd_pr__cap_mim_m3_1_C8GDQN  XC3
timestamp 0
transform 1 0 15930 0 1 -502200
box -3186 -85320 3186 85320
use sky130_fd_pr__cap_mim_m3_1_CWHDQN  XC4
timestamp 0
transform 1 0 22302 0 1 -714040
box -3186 -132720 3186 132720
use sky130_fd_pr__cap_mim_m3_1_CWHDQN  XC5
timestamp 0
transform 1 0 28674 0 1 -973280
box -3186 -132720 3186 132720
use sky130_fd_pr__cap_mim_m3_1_CWHDQN  XC6
timestamp 0
transform 1 0 35046 0 1 -1232520
box -3186 -132720 3186 132720
use sky130_fd_pr__nfet_01v8_FMMQLY  XM1
timestamp 0
transform 1 0 782 0 1 -1367886
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XM2
timestamp 0
transform 1 0 1321 0 1 -1367939
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XM3
timestamp 0
transform 1 0 1860 0 1 -1367992
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XM4
timestamp 0
transform 1 0 2399 0 1 -1368045
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XM5
timestamp 0
transform 1 0 2938 0 1 -1368098
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XM6
timestamp 0
transform 1 0 3477 0 1 -1368151
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XM7
timestamp 0
transform 1 0 4016 0 1 -1368204
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_FMMQLY  XM12
timestamp 0
transform 1 0 243 0 1 -1367833
box -296 -260 296 260
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD_1V8
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 DAC+
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 DAC-
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 I1
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 Vop
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VBP
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Von
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 VBN
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 I2
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 Clk_1
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 Clk
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 Clk_2
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 VSS
port 12 nsew
<< end >>
