*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include - Standard includes, assuming no specific fast models
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR06_main_lpe.spi
#else
.include ../../../work/xsch/CNR_GR06_main.spice
#endif

*-----------------------------------------------------------------
* OPTIONS - Operating at an elevated temperature for the fast corner
*-----------------------------------------------------------------
.option TNOM=125 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS - Defining simulation parameters, with some adjusted for fast conditions
*-----------------------------------------------------------------
.param TRF = 100p
.param t_start = 0.5u
.param t_start_del = {t_start + TRF}
.param PERIOD_CLK = 500n
.param PW_CLK = PERIOD_CLK/2

* Fast corner adjustments:
* Decreasing the threshold voltages slightly to represent faster transistor switching
.param nmos_vth_fast = 0.0   ; Adjusted for faster NMOS
.param pmos_vth_fast = -0.003 ; Adjusted for faster PMOS
.param AVDD_fast = 1.25       ; Optionally increased supply for fast corner

*-----------------------------------------------------------------
* FORCE - Applying potential fast corner conditions
*-----------------------------------------------------------------
VSS  VSS  0  dc 0
VDD  VDD_1V8 0 dc {AVDD_fast}
Vdref Vdref 0 dc 1.2

* Using adjusted threshold voltages for hypothetical signal sources (if applicable)
VT2 VT2 0 dc {nmos_vth_fast}
VT1 VT1 0 dc {pmos_vth_fast}

* Assuming other conditions remain unchanged
VBP VBP 0 dc 0.08
VBN VBN 0 dc 1.12

VCLK Clk 0 dc 0 pulse 0 1.2 {t_start} {TRF} {TRF} {PW_CLK} {PERIOD_CLK}

*-----------------------------------------------------------------
* DUT - Include the device under test as before
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE and MEASURES - Unchanged for debugging and analysis
*----------------------------------------------------------------
#ifdef Debug
.save all
#else
.save ${VPORTS}
#endif

*----------------------------------------------------------------
* NGSPICE control - Running the simulation with transient analysis
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

tran 0.1 50u 0.1u
write

run
set filetype=ascii
write "output_data_fast.txt" V(Voc)
.quit
quit

.endc

.end

