magic
tech sky130B
magscale 1 2
timestamp 1713382353
<< error_s >>
rect 2188 4783 2287 4801
rect 153 4747 2033 4783
rect 2188 4747 16283 4783
rect 79 4713 16945 4747
rect 153 4661 2033 4713
rect 2188 4679 16283 4713
rect 16415 4679 16441 4713
rect 153 4651 2044 4661
rect 147 4645 2052 4651
rect 2134 4645 16283 4679
rect 16384 4651 16441 4679
rect 16449 4661 16483 4713
rect 16615 4679 16641 4713
rect 16449 4651 16481 4661
rect 16384 4645 16481 4651
rect 143 4611 2052 4645
rect 147 4605 2052 4611
rect 153 4561 2052 4605
rect 2072 4573 2090 4577
rect 2106 4573 2124 4577
rect 2072 4561 2096 4573
rect 153 4369 2096 4561
rect 153 4325 2052 4369
rect 2072 4357 2096 4369
rect 2100 4561 2124 4573
rect 2150 4561 16283 4645
rect 16400 4611 16481 4645
rect 16600 4651 16641 4679
rect 16649 4661 16683 4713
rect 16649 4651 16681 4661
rect 16600 4645 16681 4651
rect 16791 4651 16841 4679
rect 16791 4645 16807 4651
rect 16809 4645 16877 4651
rect 16600 4611 16641 4645
rect 16649 4611 16681 4645
rect 16809 4611 16841 4645
rect 16865 4611 16875 4645
rect 16400 4605 16483 4611
rect 2100 4369 16283 4561
rect 2100 4357 2124 4369
rect 2072 4353 2090 4357
rect 2106 4353 2124 4357
rect 2150 4353 16283 4369
rect 16286 4561 16317 4577
rect 16322 4573 16327 4577
rect 16356 4573 16361 4577
rect 16366 4573 16397 4577
rect 16322 4561 16333 4573
rect 16286 4369 16333 4561
rect 16286 4353 16317 4369
rect 16322 4357 16333 4369
rect 16344 4357 16397 4573
rect 16322 4353 16327 4357
rect 16356 4353 16361 4357
rect 16366 4353 16397 4357
rect 16400 4353 16441 4605
rect 147 4319 2052 4325
rect 2134 4319 16283 4353
rect 16384 4325 16441 4353
rect 16449 4325 16483 4605
rect 16600 4605 16683 4611
rect 16486 4561 16517 4577
rect 16566 4573 16597 4577
rect 16486 4369 16527 4561
rect 16486 4353 16517 4369
rect 16529 4357 16533 4573
rect 16551 4357 16597 4573
rect 16566 4353 16597 4357
rect 16384 4319 16483 4325
rect 16600 4325 16641 4605
rect 16649 4325 16683 4605
rect 16807 4605 16877 4611
rect 16693 4353 16717 4577
rect 16773 4573 16797 4577
rect 16725 4369 16727 4561
rect 16729 4357 16733 4573
rect 16751 4357 16797 4573
rect 16773 4353 16797 4357
rect 16807 4353 16841 4605
rect 16600 4319 16683 4325
rect 16791 4325 16841 4353
rect 16791 4319 16877 4325
rect 143 4285 2052 4319
rect 147 4279 2052 4285
rect 2150 4279 16283 4319
rect 16400 4279 16481 4319
rect 16600 4285 16641 4319
rect 16649 4285 16681 4319
rect 16600 4279 16681 4285
rect 153 4269 2044 4279
rect 2152 4269 16283 4279
rect 16402 4269 16441 4279
rect 153 4217 2033 4269
rect 2188 4217 16283 4269
rect 16415 4217 16441 4269
rect 16449 4269 16481 4279
rect 16609 4269 16641 4279
rect 16449 4217 16483 4269
rect 16615 4217 16641 4269
rect 16649 4269 16681 4279
rect 16809 4285 16841 4319
rect 16865 4285 16875 4319
rect 16809 4279 16877 4285
rect 16809 4269 16841 4279
rect 16649 4217 16683 4269
rect 16830 4258 16841 4269
rect 79 4183 16945 4217
rect 153 4147 2033 4183
rect 2188 4147 16283 4183
rect 1168 3583 1274 3601
rect 4429 3583 4535 3601
rect -52 3547 1020 3583
rect 1168 3547 1834 3583
rect 2188 3547 4281 3583
rect 4429 3565 4693 3583
rect 4831 3565 15883 3583
rect 4429 3547 15952 3565
rect -52 3531 15952 3547
rect -52 3513 4701 3531
rect -52 3461 1020 3513
rect 1141 3461 1147 3513
rect 1168 3479 1852 3513
rect 1168 3461 1862 3479
rect 1984 3461 2004 3513
rect -52 3451 1091 3461
rect -52 3400 1093 3451
rect 1141 3411 1862 3461
rect 1972 3451 2004 3461
rect 2018 3479 2058 3513
rect 2188 3479 4299 3513
rect 4429 3497 4701 3513
rect 2018 3451 2068 3479
rect 2188 3461 4309 3479
rect 4429 3461 4716 3497
rect 4831 3479 15883 3531
rect 4826 3469 15883 3479
rect 2178 3451 4309 3461
rect 4419 3451 4716 3461
rect 1964 3411 2068 3451
rect 2170 3411 4309 3451
rect 4411 3429 4716 3451
rect 4823 3463 15884 3469
rect 4823 3429 15883 3463
rect 1141 3400 1852 3411
rect 1964 3405 2058 3411
rect 1964 3400 2004 3405
rect 2018 3400 2058 3405
rect 2170 3400 4299 3411
rect 4411 3400 4701 3429
rect 4823 3423 15884 3429
rect 4823 3400 15883 3423
rect -52 3377 1115 3400
rect 1119 3377 1868 3400
rect 1948 3377 2074 3400
rect 2154 3377 4315 3400
rect 4395 3395 4722 3400
rect 4802 3395 15912 3400
rect 4395 3377 4701 3395
rect -52 3361 1093 3377
rect 1141 3361 1852 3377
rect 1914 3361 1956 3373
rect 1964 3361 2004 3377
rect -52 3169 1890 3361
rect -52 3079 1093 3169
rect 1141 3153 1852 3169
rect 1892 3157 1896 3200
rect 1914 3169 2004 3361
rect 1914 3157 1956 3169
rect 1141 3085 1862 3153
rect 1964 3125 2004 3169
rect 2018 3361 2058 3377
rect 2120 3361 2162 3373
rect 2170 3361 4299 3377
rect 4361 3361 4403 3373
rect 4411 3361 4701 3377
rect 2018 3169 2096 3361
rect 2018 3153 2058 3169
rect 2098 3157 2102 3200
rect 2120 3169 4337 3361
rect 2120 3157 2162 3169
rect 2170 3153 4299 3169
rect 4339 3157 4343 3200
rect 4361 3169 4701 3361
rect 4361 3157 4403 3169
rect 4411 3153 4701 3169
rect 4709 3370 4735 3386
rect 4789 3382 4815 3386
rect 4709 3178 4744 3370
rect 4709 3162 4735 3178
rect 4746 3166 4750 3200
rect 4768 3166 4815 3382
rect 4789 3162 4815 3166
rect 2018 3125 2068 3153
rect 1964 3085 2068 3125
rect 2170 3085 4309 3153
rect 4411 3085 4716 3153
rect 4823 3125 15883 3395
rect 15899 3178 15934 3370
rect 4823 3119 15884 3125
rect 4823 3085 15883 3119
rect 1141 3079 1852 3085
rect 1964 3079 2058 3085
rect 2170 3079 4299 3085
rect 4411 3079 4701 3085
rect 4823 3079 15884 3085
rect 16013 3079 16048 3469
rect -52 3069 1091 3079
rect 1141 3069 1844 3079
rect 1972 3069 2004 3079
rect -52 3019 1020 3069
rect -52 3017 1037 3019
rect 1141 3017 1147 3069
rect 1168 3019 1852 3069
rect 1150 3017 1852 3019
rect 1984 3017 2004 3069
rect 2018 3069 2050 3079
rect 2178 3069 4291 3079
rect 4419 3069 4698 3079
rect 4826 3069 15883 3079
rect 2018 3017 2058 3069
rect 2188 3019 4299 3069
rect 4429 3019 4701 3069
rect 4831 3019 15883 3069
rect 2170 3017 4299 3019
rect 4411 3017 4701 3019
rect 4823 3017 15883 3019
rect 16013 3017 16048 3019
rect -52 2983 16048 3017
rect -52 2947 1020 2983
rect 1168 2947 1834 2983
rect 2188 2947 4281 2983
rect 4429 2947 16084 2983
rect 79 2913 16745 2947
rect 153 2861 1019 2913
rect 1158 2879 1833 2913
rect 2172 2879 4280 2913
rect 4412 2879 16083 2913
rect 16215 2879 16241 2913
rect 1125 2861 1833 2879
rect 1934 2861 1988 2879
rect 2150 2861 4280 2879
rect 153 2851 1024 2861
rect 1125 2851 1838 2861
rect 1934 2851 2044 2861
rect 2150 2851 4285 2861
rect 153 2845 1032 2851
rect 1125 2845 1846 2851
rect 1934 2845 2052 2851
rect 143 2811 1032 2845
rect 153 2801 1032 2811
rect 1141 2801 1846 2845
rect 1950 2801 2052 2845
rect 2150 2801 4293 2851
rect 4381 2845 16083 2879
rect 16184 2845 16241 2879
rect 16249 2861 16283 2913
rect 16415 2879 16441 2913
rect 16249 2845 16281 2861
rect 4397 2801 16083 2845
rect 16200 2811 16281 2845
rect 16200 2801 16241 2811
rect 63 2800 16241 2801
rect 153 2773 1032 2800
rect 1063 2773 1070 2777
rect 1097 2773 1104 2777
rect 1141 2773 1846 2800
rect 1872 2773 1884 2777
rect 1906 2773 1918 2777
rect 1950 2773 2052 2800
rect 2078 2773 2090 2777
rect 2112 2773 2124 2777
rect 2150 2773 4293 2800
rect 4319 2773 4331 2777
rect 4353 2773 4365 2777
rect 4397 2773 16083 2800
rect 16086 2773 16117 2777
rect 16122 2773 16127 2777
rect 16156 2773 16161 2777
rect 16166 2773 16197 2777
rect 16200 2773 16241 2800
rect 91 2772 137 2773
rect 153 2772 1076 2773
rect 153 2761 1032 2772
rect 1063 2761 1076 2772
rect 153 2601 1076 2761
rect 1085 2772 1890 2773
rect 1085 2761 1136 2772
rect 1141 2761 1846 2772
rect 1872 2761 1890 2772
rect 1085 2601 1890 2761
rect 1900 2772 2096 2773
rect 1900 2761 1918 2772
rect 1950 2761 2052 2772
rect 2078 2761 2096 2772
rect 1900 2601 2096 2761
rect 2106 2772 4337 2773
rect 2106 2761 2124 2772
rect 2150 2761 4293 2772
rect 4319 2761 4337 2772
rect 2106 2601 4337 2761
rect 4347 2772 16133 2773
rect 4347 2761 4365 2772
rect 4397 2761 16083 2772
rect 4347 2601 16083 2761
rect 16086 2761 16117 2772
rect 16122 2761 16133 2772
rect 16086 2601 16133 2761
rect 16144 2772 16241 2773
rect 16144 2601 16197 2772
rect 16200 2601 16241 2772
rect 16249 2801 16283 2811
rect 16400 2801 16441 2879
rect 16249 2800 16441 2801
rect 16249 2773 16283 2800
rect 16286 2773 16317 2777
rect 16366 2773 16397 2777
rect 16400 2773 16441 2800
rect 16249 2772 16333 2773
rect 16249 2601 16283 2772
rect 16286 2761 16317 2772
rect 16286 2601 16327 2761
rect 16329 2601 16333 2772
rect 16351 2772 16441 2773
rect 16351 2601 16397 2772
rect 16400 2601 16441 2772
rect 16449 2861 16483 2913
rect 16449 2811 16481 2861
rect 16591 2851 16641 2879
rect 16591 2845 16607 2851
rect 16609 2811 16641 2851
rect 16665 2811 16675 2845
rect 16449 2801 16483 2811
rect 16607 2801 16641 2811
rect 16449 2800 16641 2801
rect 16659 2800 16761 2801
rect 16449 2601 16483 2800
rect 16493 2773 16517 2777
rect 16573 2773 16597 2777
rect 16487 2772 16533 2773
rect 16493 2601 16517 2772
rect 16525 2601 16527 2761
rect 16529 2601 16533 2772
rect 16551 2772 16603 2773
rect 16551 2601 16597 2772
rect 16607 2601 16641 2800
rect 16687 2772 16733 2773
rect 16807 2601 16841 2851
rect -53 2557 16139 2601
rect 16144 2557 16841 2601
rect -53 2553 1884 2557
rect 1906 2553 2090 2557
rect 2112 2553 16083 2557
rect 16086 2553 16127 2557
rect -53 2547 1846 2553
rect 1934 2547 2052 2553
rect 2150 2547 16083 2553
rect 16147 2547 16841 2557
rect 19347 2565 19611 2583
rect 20147 2565 20411 2583
rect 19347 2547 20411 2565
rect 21547 2565 21811 2583
rect 21947 2565 22211 2583
rect 21547 2547 22211 2565
rect 23347 2565 23611 2583
rect 23747 2565 24011 2583
rect 23347 2547 24011 2565
rect 25147 2565 25411 2583
rect 25547 2565 25811 2583
rect 25147 2547 25811 2565
rect 26947 2565 27211 2583
rect 27347 2565 27611 2583
rect 26947 2547 27611 2565
rect 28747 2565 29011 2583
rect 29147 2565 29411 2583
rect 28747 2547 29411 2565
rect 30547 2565 30811 2583
rect 30947 2565 31211 2583
rect 30547 2547 31211 2565
rect 32347 2565 32611 2583
rect 32747 2565 33011 2583
rect 32347 2547 33011 2565
rect 34147 2565 34411 2583
rect 34547 2565 34811 2583
rect 34147 2547 34811 2565
rect 35947 2565 36211 2583
rect 36347 2565 36611 2583
rect 35947 2547 36611 2565
rect 37747 2565 38011 2583
rect 38147 2565 38411 2583
rect 37747 2547 38411 2565
rect 39547 2565 39811 2583
rect 39947 2565 40211 2583
rect 39547 2547 40211 2565
rect 41347 2565 41611 2583
rect 41747 2565 42011 2583
rect 41347 2547 42011 2565
rect 43147 2565 43411 2583
rect 43547 2565 43811 2583
rect 43147 2547 43811 2565
rect 44947 2565 45211 2583
rect 45347 2565 45611 2583
rect 44947 2547 45611 2565
rect 46747 2565 47011 2583
rect 47147 2565 47411 2583
rect 46747 2547 47411 2565
rect 48547 2565 48811 2583
rect 48947 2565 49211 2583
rect 48547 2547 49211 2565
rect 50347 2565 50611 2583
rect 50747 2565 51011 2583
rect 50347 2547 51011 2565
rect 52147 2565 52411 2583
rect 52547 2565 52811 2583
rect 52147 2547 52811 2565
rect 53947 2565 54211 2583
rect 54347 2565 54611 2583
rect 53947 2547 54611 2565
rect 55747 2565 56011 2583
rect 56147 2565 56411 2583
rect 55747 2547 56411 2565
rect 57547 2565 57811 2583
rect 57947 2565 58211 2583
rect 57547 2547 58211 2565
rect 59347 2565 59611 2583
rect 59747 2565 60011 2583
rect 59347 2547 60011 2565
rect 61147 2565 61411 2583
rect 61547 2565 61811 2583
rect 61147 2547 61811 2565
rect 62947 2565 63211 2583
rect 63347 2565 63611 2583
rect 62947 2547 63611 2565
rect 64747 2565 65011 2583
rect 65147 2565 65411 2583
rect 64747 2547 65411 2565
rect 66547 2565 66811 2583
rect 66947 2565 67211 2583
rect 66547 2547 67211 2565
rect 68347 2565 68611 2583
rect 68347 2547 68879 2565
rect -53 2531 68879 2547
rect -53 2513 19617 2531
rect -53 2479 1846 2513
rect 1950 2492 2052 2513
rect 2150 2492 16083 2513
rect 1941 2479 2052 2492
rect 2141 2479 16083 2492
rect 16147 2479 16841 2513
rect 16949 2479 16975 2513
rect -53 2469 1838 2479
rect 1925 2469 2044 2479
rect 2125 2469 16083 2479
rect -53 2427 1833 2469
rect 1925 2461 1983 2469
rect 2125 2461 2183 2469
rect 2188 2461 16083 2469
rect 1925 2451 2015 2461
rect 1925 2445 2017 2451
rect 2125 2445 16083 2461
rect 16125 2461 16829 2479
rect 16125 2445 16815 2461
rect 16925 2451 16975 2479
rect 16983 2461 17017 2513
rect 17149 2479 17175 2513
rect 16983 2451 17015 2461
rect 16925 2445 16941 2451
rect 16943 2445 17015 2451
rect 17125 2451 17175 2479
rect 17183 2461 17217 2513
rect 17349 2479 17375 2513
rect 17183 2451 17215 2461
rect 17125 2445 17141 2451
rect 17143 2445 17215 2451
rect 17325 2451 17375 2479
rect 17383 2461 17417 2513
rect 17549 2479 17575 2513
rect 17383 2451 17415 2461
rect 17325 2445 17341 2451
rect 17343 2445 17415 2451
rect 17525 2451 17575 2479
rect 17583 2461 17617 2513
rect 17749 2479 17775 2513
rect 17583 2451 17615 2461
rect 17525 2445 17541 2451
rect 17543 2445 17615 2451
rect 17725 2451 17775 2479
rect 17783 2461 17817 2513
rect 17949 2479 17975 2513
rect 17783 2451 17815 2461
rect 17725 2445 17741 2451
rect 17743 2445 17815 2451
rect 17925 2451 17975 2479
rect 17983 2479 18017 2513
rect 17983 2451 18033 2479
rect 18149 2461 18175 2513
rect 17925 2445 17941 2451
rect 17943 2445 18033 2451
rect 1941 2427 2017 2445
rect -53 2417 1846 2427
rect 1941 2417 2052 2427
rect 2141 2417 16083 2445
rect 16141 2417 16815 2445
rect -53 2411 16815 2417
rect 16817 2411 16841 2427
rect 16943 2411 16975 2445
rect 16983 2411 17015 2445
rect 17143 2411 17175 2445
rect 17183 2411 17215 2445
rect 17343 2411 17375 2445
rect 17383 2411 17415 2445
rect 17543 2411 17575 2445
rect 17583 2411 17615 2445
rect 17743 2411 17775 2445
rect 17783 2411 17815 2445
rect 17943 2411 17975 2445
rect 17983 2411 18033 2445
rect 18143 2451 18175 2461
rect 18183 2461 18217 2513
rect 18349 2479 18375 2513
rect 18183 2451 18215 2461
rect 18143 2445 18215 2451
rect 18325 2451 18375 2479
rect 18383 2461 18417 2513
rect 18549 2479 18575 2513
rect 18383 2451 18415 2461
rect 18325 2445 18341 2451
rect 18343 2445 18415 2451
rect 18525 2451 18575 2479
rect 18583 2461 18617 2513
rect 18749 2479 18775 2513
rect 18583 2451 18615 2461
rect 18525 2445 18541 2451
rect 18543 2445 18615 2451
rect 18725 2451 18775 2479
rect 18783 2461 18817 2513
rect 18949 2479 18975 2513
rect 18783 2451 18815 2461
rect 18725 2445 18741 2451
rect 18743 2445 18815 2451
rect 18925 2451 18975 2479
rect 18983 2461 19017 2513
rect 19149 2479 19175 2513
rect 18983 2451 19015 2461
rect 18925 2445 18941 2451
rect 18943 2445 19015 2451
rect 19125 2451 19175 2479
rect 19183 2461 19217 2513
rect 19347 2479 19617 2513
rect 19749 2497 19775 2531
rect 19183 2451 19215 2461
rect 19125 2445 19141 2451
rect 19143 2445 19215 2451
rect 19325 2451 19615 2479
rect 19725 2469 19775 2497
rect 19783 2497 19817 2531
rect 19783 2469 19833 2497
rect 19949 2479 19975 2531
rect 19725 2463 19741 2469
rect 19743 2463 19833 2469
rect 19325 2445 19341 2451
rect 18143 2411 18175 2445
rect 18183 2411 18215 2445
rect 18343 2411 18375 2445
rect 18383 2411 18415 2445
rect 18543 2411 18575 2445
rect 18583 2411 18615 2445
rect 18743 2411 18775 2445
rect 18783 2411 18815 2445
rect 18943 2411 18975 2445
rect 18983 2411 19015 2445
rect 19143 2411 19175 2445
rect 19183 2411 19215 2445
rect 19343 2420 19615 2451
rect 19743 2429 19775 2463
rect 19783 2429 19833 2463
rect 19943 2469 19975 2479
rect 19983 2479 20017 2531
rect 20147 2513 21817 2531
rect 20147 2497 20417 2513
rect 19983 2469 20015 2479
rect 19943 2463 20015 2469
rect 20125 2469 20417 2497
rect 20549 2479 20575 2513
rect 20125 2463 20141 2469
rect 19943 2429 19975 2463
rect 19983 2429 20015 2463
rect 19743 2423 19815 2429
rect 19743 2420 19775 2423
rect 19343 2411 19617 2420
rect -53 2401 16841 2411
rect 16941 2405 17017 2411
rect -53 2400 16866 2401
rect -53 2383 16841 2400
rect -53 2377 1833 2383
rect -53 2373 1861 2377
rect 1897 2373 1931 2377
rect 1941 2373 1975 2383
rect -53 2358 1873 2373
rect 1885 2358 1975 2373
rect -53 2349 1861 2358
rect -53 2347 1851 2349
rect -53 2166 531 2347
rect -53 2017 493 2166
rect 507 2162 531 2166
rect 541 2119 575 2347
rect 543 2069 575 2119
rect 549 2017 575 2069
rect 583 2119 617 2347
rect 627 2162 651 2347
rect 659 2178 661 2347
rect 663 2200 667 2347
rect 685 2166 731 2347
rect 707 2162 731 2166
rect 741 2153 775 2347
rect 725 2119 775 2153
rect 583 2069 615 2119
rect 743 2069 775 2119
rect 583 2017 617 2069
rect 749 2017 775 2069
rect 783 2153 817 2347
rect 827 2162 851 2347
rect 859 2178 861 2347
rect 863 2200 867 2347
rect 885 2166 931 2347
rect 907 2162 931 2166
rect 783 2085 833 2153
rect 941 2128 975 2347
rect 783 2069 815 2085
rect 943 2069 975 2128
rect 783 2017 817 2069
rect 949 2017 975 2069
rect 983 2128 1017 2347
rect 1027 2162 1051 2347
rect 1059 2178 1061 2347
rect 1063 2200 1067 2347
rect 1085 2166 1131 2347
rect 1107 2162 1131 2166
rect 1141 2153 1417 2347
rect 1427 2153 1451 2347
rect 1459 2169 1461 2347
rect 1463 2200 1467 2347
rect 1485 2157 1531 2347
rect 1507 2153 1531 2157
rect 1541 2153 1575 2347
rect 1125 2128 1417 2153
rect 983 2069 1015 2128
rect 1125 2119 1141 2128
rect 1143 2119 1417 2128
rect 1525 2119 1575 2153
rect 1143 2069 1415 2119
rect 1543 2069 1575 2119
rect 983 2017 1017 2069
rect 1147 2017 1417 2069
rect 1549 2017 1575 2069
rect 1583 2119 1617 2347
rect 1627 2153 1651 2347
rect 1659 2169 1661 2347
rect 1663 2200 1667 2347
rect 1685 2157 1731 2347
rect 1707 2153 1731 2157
rect 1741 2153 1775 2347
rect 1725 2119 1775 2153
rect 1583 2069 1615 2119
rect 1743 2069 1775 2119
rect 1583 2017 1617 2069
rect 1749 2017 1775 2069
rect 1783 2119 1817 2347
rect 1827 2153 1851 2347
rect 1859 2169 1861 2349
rect 1863 2200 1867 2358
rect 1885 2157 1931 2358
rect 1907 2153 1931 2157
rect 1941 2153 1975 2358
rect 1925 2119 1975 2153
rect 1783 2069 1815 2119
rect 1943 2069 1975 2119
rect 1783 2017 1817 2069
rect 1949 2017 1975 2069
rect 1983 2373 2017 2383
rect 2027 2373 2061 2377
rect 2097 2373 2131 2377
rect 2141 2373 2175 2383
rect 1983 2358 2073 2373
rect 2085 2358 2175 2373
rect 1983 2119 2017 2358
rect 2027 2349 2061 2358
rect 2027 2153 2051 2349
rect 2059 2169 2061 2349
rect 2063 2200 2067 2358
rect 2085 2157 2131 2358
rect 2107 2153 2131 2157
rect 2141 2153 2175 2358
rect 2125 2119 2175 2153
rect 1983 2069 2015 2119
rect 2143 2069 2175 2119
rect 1983 2017 2017 2069
rect 2149 2017 2175 2069
rect 2183 2347 16083 2383
rect 16097 2373 16131 2377
rect 16141 2373 16817 2383
rect 16827 2373 16861 2377
rect 16907 2373 16931 2377
rect 16085 2372 16867 2373
rect 16085 2358 16861 2372
rect 2183 2119 2217 2347
rect 2227 2153 2251 2347
rect 2259 2169 2261 2347
rect 2263 2200 2267 2347
rect 2285 2157 2331 2347
rect 2307 2153 2331 2157
rect 2341 2153 2375 2347
rect 2325 2119 2375 2153
rect 2183 2069 2215 2119
rect 2343 2069 2375 2119
rect 2183 2017 2217 2069
rect 2349 2017 2375 2069
rect 2383 2119 2417 2347
rect 2427 2153 2451 2347
rect 2459 2169 2461 2347
rect 2463 2200 2467 2347
rect 2485 2157 2531 2347
rect 2507 2153 2531 2157
rect 2541 2153 2575 2347
rect 2525 2119 2575 2153
rect 2383 2069 2415 2119
rect 2543 2069 2575 2119
rect 2383 2017 2417 2069
rect 2549 2017 2575 2069
rect 2583 2153 2617 2347
rect 2627 2153 2651 2347
rect 2659 2169 2661 2347
rect 2663 2200 2667 2347
rect 2685 2157 2731 2347
rect 2707 2153 2731 2157
rect 2583 2085 2633 2153
rect 2741 2119 2775 2347
rect 2583 2069 2615 2085
rect 2743 2069 2775 2119
rect 2583 2017 2617 2069
rect 2749 2017 2775 2069
rect 2783 2119 2817 2347
rect 2827 2153 2851 2347
rect 2859 2169 2861 2347
rect 2863 2200 2867 2347
rect 2885 2157 2931 2347
rect 2907 2153 2931 2157
rect 2941 2153 2975 2347
rect 2925 2119 2975 2153
rect 2783 2069 2815 2119
rect 2943 2069 2975 2119
rect 2783 2017 2817 2069
rect 2949 2017 2975 2069
rect 2983 2119 3017 2347
rect 3027 2153 3051 2347
rect 3059 2169 3061 2347
rect 3063 2200 3067 2347
rect 3085 2157 3131 2347
rect 3107 2153 3131 2157
rect 3141 2153 3175 2347
rect 3125 2119 3175 2153
rect 2983 2069 3015 2119
rect 3143 2069 3175 2119
rect 2983 2017 3017 2069
rect 3149 2017 3175 2069
rect 3183 2119 3217 2347
rect 3227 2153 3251 2347
rect 3259 2169 3261 2347
rect 3263 2200 3267 2347
rect 3285 2157 3331 2347
rect 3307 2153 3331 2157
rect 3341 2153 3375 2347
rect 3325 2119 3375 2153
rect 3183 2069 3215 2119
rect 3343 2069 3375 2119
rect 3183 2017 3217 2069
rect 3349 2017 3375 2069
rect 3383 2119 3417 2347
rect 3427 2153 3451 2347
rect 3459 2169 3461 2347
rect 3463 2200 3467 2347
rect 3485 2157 3531 2347
rect 3507 2153 3531 2157
rect 3541 2153 3575 2347
rect 3525 2119 3575 2153
rect 3383 2069 3415 2119
rect 3543 2069 3575 2119
rect 3383 2017 3417 2069
rect 3549 2017 3575 2069
rect 3583 2119 3617 2347
rect 3627 2153 3651 2347
rect 3659 2169 3661 2347
rect 3663 2200 3667 2347
rect 3685 2157 3731 2347
rect 3707 2153 3731 2157
rect 3741 2153 3775 2347
rect 3725 2119 3775 2153
rect 3583 2069 3615 2119
rect 3743 2069 3775 2119
rect 3583 2017 3617 2069
rect 3749 2017 3775 2069
rect 3783 2119 3817 2347
rect 3827 2153 3851 2347
rect 3859 2169 3861 2347
rect 3863 2200 3867 2347
rect 3885 2157 3931 2347
rect 3907 2153 3931 2157
rect 3941 2153 4217 2347
rect 4227 2162 4251 2347
rect 4259 2178 4261 2347
rect 4263 2200 4267 2347
rect 4285 2166 4331 2347
rect 4307 2162 4331 2166
rect 4341 2153 4375 2347
rect 3925 2128 4217 2153
rect 4325 2128 4375 2153
rect 3925 2119 4215 2128
rect 4325 2119 4341 2128
rect 3783 2069 3815 2119
rect 3943 2069 4215 2119
rect 4343 2069 4375 2128
rect 3783 2017 3817 2069
rect 3947 2017 4217 2069
rect 4349 2017 4375 2069
rect 4383 2153 4417 2347
rect 4427 2162 4451 2347
rect 4459 2178 4461 2347
rect 4463 2200 4467 2347
rect 4485 2166 4531 2347
rect 4507 2162 4531 2166
rect 4383 2085 4433 2153
rect 4541 2119 4575 2347
rect 4383 2069 4415 2085
rect 4543 2069 4575 2119
rect 4383 2017 4417 2069
rect 4549 2017 4575 2069
rect 4583 2119 4617 2347
rect 4627 2162 4651 2347
rect 4659 2178 4661 2347
rect 4663 2200 4667 2347
rect 4685 2166 4731 2347
rect 4707 2162 4731 2166
rect 4741 2153 5017 2347
rect 5027 2153 5051 2347
rect 5059 2169 5061 2347
rect 5063 2200 5067 2347
rect 5085 2157 5131 2347
rect 5107 2153 5131 2157
rect 5141 2153 5175 2347
rect 4725 2119 5017 2153
rect 5125 2119 5175 2153
rect 4583 2069 4615 2119
rect 4743 2069 5015 2119
rect 5143 2069 5175 2119
rect 4583 2017 4617 2069
rect 4747 2017 5017 2069
rect 5149 2017 5175 2069
rect 5183 2119 5217 2347
rect 5227 2153 5251 2347
rect 5259 2169 5261 2347
rect 5263 2200 5267 2347
rect 5285 2157 5331 2347
rect 5307 2153 5331 2157
rect 5341 2153 5375 2347
rect 5325 2119 5375 2153
rect 5183 2069 5215 2119
rect 5343 2069 5375 2119
rect 5183 2017 5217 2069
rect 5349 2017 5375 2069
rect 5383 2119 5417 2347
rect 5427 2153 5451 2347
rect 5459 2169 5461 2347
rect 5463 2200 5467 2347
rect 5485 2157 5531 2347
rect 5507 2153 5531 2157
rect 5541 2153 5575 2347
rect 5525 2119 5575 2153
rect 5383 2069 5415 2119
rect 5543 2069 5575 2119
rect 5383 2017 5417 2069
rect 5549 2017 5575 2069
rect 5583 2119 5617 2347
rect 5627 2153 5651 2347
rect 5659 2169 5661 2347
rect 5663 2200 5667 2347
rect 5685 2157 5731 2347
rect 5707 2153 5731 2157
rect 5741 2153 5775 2347
rect 5725 2119 5775 2153
rect 5583 2069 5615 2119
rect 5743 2069 5775 2119
rect 5583 2017 5617 2069
rect 5749 2017 5775 2069
rect 5783 2119 5817 2347
rect 5827 2153 5851 2347
rect 5859 2169 5861 2347
rect 5863 2200 5867 2347
rect 5885 2157 5931 2347
rect 5907 2153 5931 2157
rect 5941 2153 5975 2347
rect 5925 2119 5975 2153
rect 5783 2069 5815 2119
rect 5943 2069 5975 2119
rect 5783 2017 5817 2069
rect 5949 2017 5975 2069
rect 5983 2119 6017 2347
rect 6027 2153 6051 2347
rect 6059 2169 6061 2347
rect 6063 2200 6067 2347
rect 6085 2157 6131 2347
rect 6107 2153 6131 2157
rect 6141 2153 6175 2347
rect 6125 2119 6175 2153
rect 5983 2069 6015 2119
rect 6143 2069 6175 2119
rect 5983 2017 6017 2069
rect 6149 2017 6175 2069
rect 6183 2153 6217 2347
rect 6227 2153 6251 2347
rect 6259 2169 6261 2347
rect 6263 2200 6267 2347
rect 6285 2157 6331 2347
rect 6307 2153 6331 2157
rect 6183 2085 6233 2153
rect 6341 2119 6375 2347
rect 6183 2069 6215 2085
rect 6343 2069 6375 2119
rect 6183 2017 6217 2069
rect 6349 2017 6375 2069
rect 6383 2119 6417 2347
rect 6427 2153 6451 2347
rect 6459 2169 6461 2347
rect 6463 2200 6467 2347
rect 6485 2157 6531 2347
rect 6507 2153 6531 2157
rect 6541 2153 6575 2347
rect 6525 2119 6575 2153
rect 6383 2069 6415 2119
rect 6543 2069 6575 2119
rect 6383 2017 6417 2069
rect 6549 2017 6575 2069
rect 6583 2119 6617 2347
rect 6627 2153 6651 2347
rect 6659 2169 6661 2347
rect 6663 2200 6667 2347
rect 6685 2157 6731 2347
rect 6707 2153 6731 2157
rect 6741 2153 6775 2347
rect 6725 2119 6775 2153
rect 6583 2069 6615 2119
rect 6743 2069 6775 2119
rect 6583 2017 6617 2069
rect 6749 2017 6775 2069
rect 6783 2119 6817 2347
rect 6827 2153 6851 2347
rect 6859 2169 6861 2347
rect 6863 2200 6867 2347
rect 6885 2157 6931 2347
rect 6907 2153 6931 2157
rect 6941 2153 6975 2347
rect 6925 2119 6975 2153
rect 6783 2069 6815 2119
rect 6943 2069 6975 2119
rect 6783 2017 6817 2069
rect 6949 2017 6975 2069
rect 6983 2119 7017 2347
rect 7027 2153 7051 2347
rect 7059 2169 7061 2347
rect 7063 2200 7067 2347
rect 7085 2157 7131 2347
rect 7107 2153 7131 2157
rect 7141 2153 7175 2347
rect 7125 2119 7175 2153
rect 6983 2069 7015 2119
rect 7143 2069 7175 2119
rect 6983 2017 7017 2069
rect 7149 2017 7175 2069
rect 7183 2119 7217 2347
rect 7227 2153 7251 2347
rect 7259 2169 7261 2347
rect 7263 2200 7267 2347
rect 7285 2157 7331 2347
rect 7307 2153 7331 2157
rect 7341 2153 7375 2347
rect 7325 2119 7375 2153
rect 7183 2069 7215 2119
rect 7343 2069 7375 2119
rect 7183 2017 7217 2069
rect 7349 2017 7375 2069
rect 7383 2119 7417 2347
rect 7427 2153 7451 2347
rect 7459 2169 7461 2347
rect 7463 2200 7467 2347
rect 7485 2157 7531 2347
rect 7507 2153 7531 2157
rect 7541 2153 7575 2347
rect 7525 2119 7575 2153
rect 7383 2069 7415 2119
rect 7543 2069 7575 2119
rect 7383 2017 7417 2069
rect 7549 2017 7575 2069
rect 7583 2153 7617 2347
rect 7627 2153 7651 2347
rect 7659 2169 7661 2347
rect 7663 2200 7667 2347
rect 7685 2157 7731 2347
rect 7707 2153 7731 2157
rect 7583 2085 7633 2153
rect 7741 2119 7775 2347
rect 7583 2069 7615 2085
rect 7743 2069 7775 2119
rect 7583 2017 7617 2069
rect 7749 2017 7775 2069
rect 7783 2119 7817 2347
rect 7827 2153 7851 2347
rect 7859 2169 7861 2347
rect 7863 2200 7867 2347
rect 7885 2157 7931 2347
rect 7907 2153 7931 2157
rect 7941 2153 7975 2347
rect 7925 2119 7975 2153
rect 7783 2069 7815 2119
rect 7943 2069 7975 2119
rect 7783 2017 7817 2069
rect 7949 2017 7975 2069
rect 7983 2119 8017 2347
rect 8027 2153 8051 2347
rect 8059 2169 8061 2347
rect 8063 2200 8067 2347
rect 8085 2157 8131 2347
rect 8107 2153 8131 2157
rect 8141 2153 8175 2347
rect 8125 2119 8175 2153
rect 7983 2069 8015 2119
rect 8143 2069 8175 2119
rect 7983 2017 8017 2069
rect 8149 2017 8175 2069
rect 8183 2119 8217 2347
rect 8227 2153 8251 2347
rect 8259 2169 8261 2347
rect 8263 2200 8267 2347
rect 8285 2157 8331 2347
rect 8307 2153 8331 2157
rect 8341 2153 8375 2347
rect 8325 2119 8375 2153
rect 8183 2069 8215 2119
rect 8343 2069 8375 2119
rect 8183 2017 8217 2069
rect 8349 2017 8375 2069
rect 8383 2119 8417 2347
rect 8427 2153 8451 2347
rect 8459 2169 8461 2347
rect 8463 2200 8467 2347
rect 8485 2157 8531 2347
rect 8507 2153 8531 2157
rect 8541 2153 8575 2347
rect 8525 2119 8575 2153
rect 8383 2069 8415 2119
rect 8543 2069 8575 2119
rect 8383 2017 8417 2069
rect 8549 2017 8575 2069
rect 8583 2119 8617 2347
rect 8627 2153 8651 2347
rect 8659 2169 8661 2347
rect 8663 2200 8667 2347
rect 8685 2157 8731 2347
rect 8707 2153 8731 2157
rect 8741 2153 8775 2347
rect 8725 2119 8775 2153
rect 8583 2069 8615 2119
rect 8743 2069 8775 2119
rect 8583 2017 8617 2069
rect 8749 2017 8775 2069
rect 8783 2119 8817 2347
rect 8827 2153 8851 2347
rect 8859 2169 8861 2347
rect 8863 2200 8867 2347
rect 8885 2157 8931 2347
rect 8907 2153 8931 2157
rect 8941 2153 9217 2347
rect 9227 2162 9251 2347
rect 9259 2178 9261 2347
rect 9263 2200 9267 2347
rect 9285 2166 9331 2347
rect 9307 2162 9331 2166
rect 9341 2153 9617 2347
rect 9627 2153 9651 2347
rect 9659 2169 9661 2347
rect 9663 2200 9667 2347
rect 9685 2157 9731 2347
rect 9707 2153 9731 2157
rect 9741 2153 9775 2347
rect 8925 2128 9217 2153
rect 8925 2119 9215 2128
rect 9325 2119 9617 2153
rect 9725 2119 9775 2153
rect 8783 2069 8815 2119
rect 8943 2069 9215 2119
rect 9343 2069 9615 2119
rect 9743 2069 9775 2119
rect 8783 2017 8817 2069
rect 8947 2017 9217 2069
rect 9347 2017 9617 2069
rect 9749 2017 9775 2069
rect 9783 2119 9817 2347
rect 9827 2153 9851 2347
rect 9859 2169 9861 2347
rect 9863 2200 9867 2347
rect 9885 2157 9931 2347
rect 9907 2153 9931 2157
rect 9941 2153 9975 2347
rect 9925 2119 9975 2153
rect 9783 2069 9815 2119
rect 9943 2069 9975 2119
rect 9783 2017 9817 2069
rect 9949 2017 9975 2069
rect 9983 2119 10017 2347
rect 10027 2153 10051 2347
rect 10059 2169 10061 2347
rect 10063 2200 10067 2347
rect 10085 2157 10131 2347
rect 10107 2153 10131 2157
rect 10141 2153 10175 2347
rect 10125 2119 10175 2153
rect 9983 2069 10015 2119
rect 10143 2069 10175 2119
rect 9983 2017 10017 2069
rect 10149 2017 10175 2069
rect 10183 2119 10217 2347
rect 10227 2153 10251 2347
rect 10259 2169 10261 2347
rect 10263 2200 10267 2347
rect 10285 2157 10331 2347
rect 10307 2153 10331 2157
rect 10341 2153 10375 2347
rect 10325 2119 10375 2153
rect 10183 2069 10215 2119
rect 10343 2069 10375 2119
rect 10183 2017 10217 2069
rect 10349 2017 10375 2069
rect 10383 2119 10417 2347
rect 10427 2153 10451 2347
rect 10459 2169 10461 2347
rect 10463 2200 10467 2347
rect 10485 2157 10531 2347
rect 10507 2153 10531 2157
rect 10541 2153 10575 2347
rect 10525 2119 10575 2153
rect 10383 2069 10415 2119
rect 10543 2069 10575 2119
rect 10383 2017 10417 2069
rect 10549 2017 10575 2069
rect 10583 2119 10617 2347
rect 10627 2153 10651 2347
rect 10659 2169 10661 2347
rect 10663 2200 10667 2347
rect 10685 2157 10731 2347
rect 10707 2153 10731 2157
rect 10741 2153 11017 2347
rect 11027 2162 11051 2347
rect 11059 2178 11061 2347
rect 11063 2200 11067 2347
rect 11085 2166 11131 2347
rect 11107 2162 11131 2166
rect 11141 2153 11417 2347
rect 11427 2153 11451 2347
rect 11459 2169 11461 2347
rect 11463 2200 11467 2347
rect 11485 2157 11531 2347
rect 11507 2153 11531 2157
rect 11541 2153 11575 2347
rect 10725 2119 11017 2153
rect 11125 2128 11417 2153
rect 11125 2119 11141 2128
rect 11143 2119 11417 2128
rect 11525 2119 11575 2153
rect 10583 2069 10615 2119
rect 10743 2069 11015 2119
rect 11143 2069 11415 2119
rect 11543 2069 11575 2119
rect 10583 2017 10617 2069
rect 10747 2017 11017 2069
rect 11147 2017 11417 2069
rect 11549 2017 11575 2069
rect 11583 2119 11617 2347
rect 11627 2153 11651 2347
rect 11659 2169 11661 2347
rect 11663 2200 11667 2347
rect 11685 2157 11731 2347
rect 11707 2153 11731 2157
rect 11741 2153 11775 2347
rect 11725 2119 11775 2153
rect 11583 2069 11615 2119
rect 11743 2069 11775 2119
rect 11583 2017 11617 2069
rect 11749 2017 11775 2069
rect 11783 2119 11817 2347
rect 11827 2153 11851 2347
rect 11859 2169 11861 2347
rect 11863 2200 11867 2347
rect 11885 2157 11931 2347
rect 11907 2153 11931 2157
rect 11941 2153 11975 2347
rect 11925 2119 11975 2153
rect 11783 2069 11815 2119
rect 11943 2069 11975 2119
rect 11783 2017 11817 2069
rect 11949 2017 11975 2069
rect 11983 2119 12017 2347
rect 12027 2153 12051 2347
rect 12059 2169 12061 2347
rect 12063 2200 12067 2347
rect 12085 2157 12131 2347
rect 12107 2153 12131 2157
rect 12141 2153 12175 2347
rect 12125 2119 12175 2153
rect 11983 2069 12015 2119
rect 12143 2069 12175 2119
rect 11983 2017 12017 2069
rect 12149 2017 12175 2069
rect 12183 2119 12217 2347
rect 12227 2153 12251 2347
rect 12259 2169 12261 2347
rect 12263 2200 12267 2347
rect 12285 2157 12331 2347
rect 12307 2153 12331 2157
rect 12341 2153 12375 2347
rect 12325 2119 12375 2153
rect 12183 2069 12215 2119
rect 12343 2069 12375 2119
rect 12183 2017 12217 2069
rect 12349 2017 12375 2069
rect 12383 2119 12417 2347
rect 12427 2153 12451 2347
rect 12459 2169 12461 2347
rect 12463 2200 12467 2347
rect 12485 2157 12531 2347
rect 12507 2153 12531 2157
rect 12541 2153 12817 2347
rect 12827 2162 12851 2347
rect 12859 2178 12861 2347
rect 12863 2200 12867 2347
rect 12885 2166 12931 2347
rect 12907 2162 12931 2166
rect 12941 2153 13217 2347
rect 13227 2153 13251 2347
rect 13259 2169 13261 2347
rect 13263 2200 13267 2347
rect 13285 2157 13331 2347
rect 13307 2153 13331 2157
rect 13341 2153 13375 2347
rect 12525 2128 12817 2153
rect 12525 2119 12815 2128
rect 12925 2119 13217 2153
rect 13325 2119 13375 2153
rect 12383 2069 12415 2119
rect 12543 2069 12815 2119
rect 12943 2069 13215 2119
rect 13343 2069 13375 2119
rect 12383 2017 12417 2069
rect 12547 2017 12817 2069
rect 12947 2017 13217 2069
rect 13349 2017 13375 2069
rect 13383 2119 13417 2347
rect 13427 2153 13451 2347
rect 13459 2169 13461 2347
rect 13463 2200 13467 2347
rect 13485 2157 13531 2347
rect 13507 2153 13531 2157
rect 13541 2153 13575 2347
rect 13525 2119 13575 2153
rect 13383 2069 13415 2119
rect 13543 2069 13575 2119
rect 13383 2017 13417 2069
rect 13549 2017 13575 2069
rect 13583 2119 13617 2347
rect 13627 2153 13651 2347
rect 13659 2169 13661 2347
rect 13663 2200 13667 2347
rect 13685 2157 13731 2347
rect 13707 2153 13731 2157
rect 13741 2153 13775 2347
rect 13725 2119 13775 2153
rect 13583 2069 13615 2119
rect 13743 2069 13775 2119
rect 13583 2017 13617 2069
rect 13749 2017 13775 2069
rect 13783 2119 13817 2347
rect 13827 2153 13851 2347
rect 13859 2169 13861 2347
rect 13863 2200 13867 2347
rect 13885 2157 13931 2347
rect 13907 2153 13931 2157
rect 13941 2153 13975 2347
rect 13925 2119 13975 2153
rect 13783 2069 13815 2119
rect 13943 2069 13975 2119
rect 13783 2017 13817 2069
rect 13949 2017 13975 2069
rect 13983 2119 14017 2347
rect 14027 2153 14051 2347
rect 14059 2169 14061 2347
rect 14063 2200 14067 2347
rect 14085 2157 14131 2347
rect 14107 2153 14131 2157
rect 14141 2153 14175 2347
rect 14125 2119 14175 2153
rect 13983 2069 14015 2119
rect 14143 2069 14175 2119
rect 13983 2017 14017 2069
rect 14149 2017 14175 2069
rect 14183 2119 14217 2347
rect 14227 2153 14251 2347
rect 14259 2169 14261 2347
rect 14263 2200 14267 2347
rect 14285 2157 14331 2347
rect 14307 2153 14331 2157
rect 14341 2153 14617 2347
rect 14627 2162 14651 2347
rect 14659 2178 14661 2347
rect 14663 2200 14667 2347
rect 14685 2166 14731 2347
rect 14707 2162 14731 2166
rect 14741 2153 15017 2347
rect 15027 2153 15051 2347
rect 15059 2169 15061 2347
rect 15063 2200 15067 2347
rect 15085 2157 15131 2347
rect 15107 2153 15131 2157
rect 15141 2153 15175 2347
rect 14325 2119 14617 2153
rect 14725 2128 15017 2153
rect 14725 2119 14741 2128
rect 14743 2119 15017 2128
rect 15125 2119 15175 2153
rect 14183 2069 14215 2119
rect 14343 2069 14615 2119
rect 14743 2069 15015 2119
rect 15143 2069 15175 2119
rect 14183 2017 14217 2069
rect 14347 2017 14617 2069
rect 14747 2017 15017 2069
rect 15149 2017 15175 2069
rect 15183 2119 15217 2347
rect 15227 2153 15251 2347
rect 15259 2169 15261 2347
rect 15263 2200 15267 2347
rect 15285 2157 15331 2347
rect 15307 2153 15331 2157
rect 15341 2153 15375 2347
rect 15325 2119 15375 2153
rect 15183 2069 15215 2119
rect 15343 2069 15375 2119
rect 15183 2017 15217 2069
rect 15349 2017 15375 2069
rect 15383 2119 15417 2347
rect 15427 2153 15451 2347
rect 15459 2169 15461 2347
rect 15463 2200 15467 2347
rect 15485 2157 15531 2347
rect 15507 2153 15531 2157
rect 15541 2153 15575 2347
rect 15525 2119 15575 2153
rect 15383 2069 15415 2119
rect 15543 2069 15575 2119
rect 15383 2017 15417 2069
rect 15549 2017 15575 2069
rect 15583 2119 15617 2347
rect 15627 2153 15651 2347
rect 15659 2169 15661 2347
rect 15663 2200 15667 2347
rect 15685 2157 15731 2347
rect 15707 2153 15731 2157
rect 15741 2153 15775 2347
rect 15725 2119 15775 2153
rect 15583 2069 15615 2119
rect 15743 2069 15775 2119
rect 15583 2017 15617 2069
rect 15749 2017 15775 2069
rect 15783 2119 15817 2347
rect 15827 2153 15851 2347
rect 15859 2169 15861 2347
rect 15863 2200 15867 2347
rect 15863 2129 15873 2200
rect 15885 2157 15931 2347
rect 15907 2153 15931 2157
rect 15941 2153 15975 2347
rect 15925 2125 15975 2153
rect 15983 2125 16017 2347
rect 16027 2153 16051 2347
rect 16059 2169 16061 2347
rect 16063 2157 16067 2347
rect 16085 2157 16131 2358
rect 16107 2153 16131 2157
rect 16141 2347 16817 2358
rect 16141 2153 16417 2347
rect 16427 2162 16451 2347
rect 16459 2178 16461 2347
rect 16463 2166 16467 2347
rect 16485 2166 16531 2347
rect 16507 2162 16531 2166
rect 16541 2153 16817 2347
rect 16827 2349 16861 2358
rect 16827 2153 16851 2349
rect 16859 2169 16861 2349
rect 16863 2157 16867 2372
rect 16885 2157 16931 2373
rect 16907 2153 16931 2157
rect 16941 2153 16975 2405
rect 15925 2119 16017 2125
rect 16125 2128 16417 2153
rect 16525 2128 16817 2153
rect 16125 2119 16415 2128
rect 16525 2119 16541 2128
rect 16543 2119 16817 2128
rect 16925 2125 16975 2153
rect 16983 2125 17017 2405
rect 17141 2405 17217 2411
rect 17027 2153 17051 2377
rect 17107 2373 17131 2377
rect 17059 2169 17061 2361
rect 17063 2157 17067 2373
rect 17085 2157 17131 2373
rect 17107 2153 17131 2157
rect 17141 2153 17175 2405
rect 16925 2119 17017 2125
rect 17125 2125 17175 2153
rect 17183 2125 17217 2405
rect 17341 2405 17417 2411
rect 17227 2153 17251 2377
rect 17307 2373 17331 2377
rect 17259 2169 17261 2361
rect 17263 2157 17267 2373
rect 17285 2157 17331 2373
rect 17307 2153 17331 2157
rect 17341 2153 17375 2405
rect 17125 2119 17217 2125
rect 17325 2125 17375 2153
rect 17383 2125 17417 2405
rect 17541 2405 17617 2411
rect 17427 2153 17451 2377
rect 17507 2373 17531 2377
rect 17459 2169 17461 2361
rect 17463 2157 17467 2373
rect 17485 2157 17531 2373
rect 17507 2153 17531 2157
rect 17541 2153 17575 2405
rect 17325 2119 17417 2125
rect 17525 2125 17575 2153
rect 17583 2125 17617 2405
rect 17741 2405 17817 2411
rect 17627 2153 17651 2377
rect 17707 2373 17731 2377
rect 17659 2169 17661 2361
rect 17663 2157 17667 2373
rect 17685 2157 17731 2373
rect 17707 2153 17731 2157
rect 17741 2153 17775 2405
rect 17525 2119 17617 2125
rect 17725 2125 17775 2153
rect 17783 2125 17817 2405
rect 17941 2405 18017 2411
rect 17827 2153 17851 2377
rect 17907 2373 17931 2377
rect 17859 2169 17861 2361
rect 17863 2157 17867 2373
rect 17885 2157 17931 2373
rect 17907 2153 17931 2157
rect 17941 2153 17975 2405
rect 17725 2119 17817 2125
rect 17925 2125 17975 2153
rect 17983 2153 18017 2405
rect 18141 2405 18217 2411
rect 18027 2153 18051 2377
rect 18107 2373 18131 2377
rect 18059 2169 18061 2361
rect 18063 2157 18067 2373
rect 18085 2157 18131 2373
rect 18107 2153 18131 2157
rect 17983 2125 18033 2153
rect 17925 2119 18033 2125
rect 18141 2125 18175 2405
rect 18183 2125 18217 2405
rect 18341 2405 18417 2411
rect 18227 2153 18251 2377
rect 18307 2373 18331 2377
rect 18259 2169 18261 2361
rect 18263 2157 18267 2373
rect 18285 2157 18331 2373
rect 18307 2153 18331 2157
rect 18341 2153 18375 2405
rect 18141 2119 18217 2125
rect 18325 2125 18375 2153
rect 18383 2125 18417 2405
rect 18541 2405 18617 2411
rect 18427 2153 18451 2377
rect 18507 2373 18531 2377
rect 18459 2169 18461 2361
rect 18463 2157 18467 2373
rect 18485 2157 18531 2373
rect 18507 2153 18531 2157
rect 18541 2153 18575 2405
rect 18325 2119 18417 2125
rect 18525 2125 18575 2153
rect 18583 2125 18617 2405
rect 18741 2405 18817 2411
rect 18627 2153 18651 2377
rect 18707 2373 18731 2377
rect 18659 2169 18661 2361
rect 18663 2157 18667 2373
rect 18685 2157 18731 2373
rect 18707 2153 18731 2157
rect 18741 2153 18775 2405
rect 18525 2119 18617 2125
rect 18725 2125 18775 2153
rect 18783 2125 18817 2405
rect 18941 2405 19017 2411
rect 18827 2153 18851 2377
rect 18907 2373 18931 2377
rect 18859 2169 18861 2361
rect 18863 2157 18867 2373
rect 18885 2157 18931 2373
rect 18907 2153 18931 2157
rect 18941 2153 18975 2405
rect 18725 2119 18817 2125
rect 18925 2125 18975 2153
rect 18983 2125 19017 2405
rect 19141 2405 19217 2411
rect 19027 2153 19051 2377
rect 19107 2373 19131 2377
rect 19059 2169 19061 2361
rect 19063 2157 19067 2373
rect 19085 2157 19131 2373
rect 19107 2153 19131 2157
rect 19141 2153 19175 2405
rect 18925 2119 19017 2125
rect 19125 2125 19175 2153
rect 19183 2125 19217 2405
rect 19227 2153 19251 2377
rect 19307 2373 19331 2377
rect 19259 2169 19261 2361
rect 19263 2157 19267 2373
rect 19285 2157 19331 2373
rect 19307 2153 19331 2157
rect 19341 2153 19617 2411
rect 19627 2162 19651 2386
rect 19707 2382 19731 2386
rect 19659 2178 19661 2370
rect 19663 2166 19667 2382
rect 19685 2166 19731 2382
rect 19707 2162 19731 2166
rect 19741 2153 19775 2420
rect 19125 2119 19217 2125
rect 19325 2128 19617 2153
rect 19725 2128 19775 2153
rect 19325 2119 19615 2128
rect 19725 2119 19741 2128
rect 19743 2125 19775 2128
rect 19783 2420 19815 2423
rect 19943 2423 20015 2429
rect 19943 2420 19975 2423
rect 19783 2153 19817 2420
rect 19827 2162 19851 2386
rect 19907 2382 19931 2386
rect 19859 2178 19861 2370
rect 19863 2166 19867 2382
rect 19885 2166 19931 2382
rect 19907 2162 19931 2166
rect 19783 2125 19833 2153
rect 19941 2128 19975 2420
rect 19743 2119 19833 2125
rect 15783 2069 15815 2119
rect 15943 2085 15975 2119
rect 15983 2085 16015 2119
rect 15943 2079 16015 2085
rect 15943 2069 15975 2079
rect 15783 2017 15817 2069
rect 15949 2017 15975 2069
rect 15983 2069 16015 2079
rect 16143 2069 16415 2119
rect 16543 2069 16815 2119
rect 16943 2085 16975 2119
rect 16983 2085 17015 2119
rect 16943 2079 17015 2085
rect 16943 2069 16975 2079
rect 15983 2017 16017 2069
rect 16147 2017 16417 2069
rect 16547 2017 16817 2069
rect 16949 2017 16975 2069
rect 16983 2069 17015 2079
rect 17143 2085 17175 2119
rect 17183 2085 17215 2119
rect 17143 2079 17215 2085
rect 17143 2069 17175 2079
rect 16983 2017 17017 2069
rect 17149 2017 17175 2069
rect 17183 2069 17215 2079
rect 17343 2085 17375 2119
rect 17383 2085 17415 2119
rect 17343 2079 17415 2085
rect 17343 2069 17375 2079
rect 17183 2017 17217 2069
rect 17349 2017 17375 2069
rect 17383 2069 17415 2079
rect 17543 2085 17575 2119
rect 17583 2085 17615 2119
rect 17543 2079 17615 2085
rect 17543 2069 17575 2079
rect 17383 2017 17417 2069
rect 17549 2017 17575 2069
rect 17583 2069 17615 2079
rect 17743 2085 17775 2119
rect 17783 2085 17815 2119
rect 17743 2079 17815 2085
rect 17743 2069 17775 2079
rect 17583 2017 17617 2069
rect 17749 2017 17775 2069
rect 17783 2069 17815 2079
rect 17943 2085 17975 2119
rect 17983 2085 18033 2119
rect 18143 2085 18175 2119
rect 18183 2085 18215 2119
rect 17943 2079 18015 2085
rect 17943 2069 17975 2079
rect 17783 2017 17817 2069
rect 17949 2017 17975 2069
rect 17983 2069 18015 2079
rect 18143 2079 18215 2085
rect 18143 2069 18175 2079
rect 17983 2017 18017 2069
rect 18149 2017 18175 2069
rect 18183 2069 18215 2079
rect 18343 2085 18375 2119
rect 18383 2085 18415 2119
rect 18343 2079 18415 2085
rect 18343 2069 18375 2079
rect 18183 2017 18217 2069
rect 18349 2017 18375 2069
rect 18383 2069 18415 2079
rect 18543 2085 18575 2119
rect 18583 2085 18615 2119
rect 18543 2079 18615 2085
rect 18543 2069 18575 2079
rect 18383 2017 18417 2069
rect 18549 2017 18575 2069
rect 18583 2069 18615 2079
rect 18743 2085 18775 2119
rect 18783 2085 18815 2119
rect 18743 2079 18815 2085
rect 18743 2069 18775 2079
rect 18583 2017 18617 2069
rect 18749 2017 18775 2069
rect 18783 2069 18815 2079
rect 18943 2085 18975 2119
rect 18983 2085 19015 2119
rect 18943 2079 19015 2085
rect 18943 2069 18975 2079
rect 18783 2017 18817 2069
rect 18949 2017 18975 2069
rect 18983 2069 19015 2079
rect 19143 2085 19175 2119
rect 19183 2085 19215 2119
rect 19143 2079 19215 2085
rect 19143 2069 19175 2079
rect 18983 2017 19017 2069
rect 19149 2017 19175 2069
rect 19183 2069 19215 2079
rect 19343 2069 19615 2119
rect 19743 2085 19775 2119
rect 19783 2085 19833 2119
rect 19943 2125 19975 2128
rect 19983 2420 20015 2423
rect 20143 2461 20417 2469
rect 20143 2420 20415 2461
rect 20525 2451 20575 2479
rect 20583 2461 20617 2513
rect 20749 2479 20775 2513
rect 20583 2451 20615 2461
rect 20525 2445 20541 2451
rect 20543 2445 20615 2451
rect 20725 2451 20775 2479
rect 20783 2461 20817 2513
rect 20949 2479 20975 2513
rect 20783 2451 20815 2461
rect 20725 2445 20741 2451
rect 20743 2445 20815 2451
rect 20925 2451 20975 2479
rect 20983 2461 21017 2513
rect 21149 2479 21175 2513
rect 20983 2451 21015 2461
rect 20925 2445 20941 2451
rect 20943 2445 21015 2451
rect 21125 2451 21175 2479
rect 21183 2461 21217 2513
rect 21349 2479 21375 2513
rect 21183 2451 21215 2461
rect 21125 2445 21141 2451
rect 21143 2445 21215 2451
rect 21325 2451 21375 2479
rect 21383 2461 21417 2513
rect 21547 2479 21817 2513
rect 21947 2513 23617 2531
rect 21947 2497 22217 2513
rect 21383 2451 21415 2461
rect 21325 2445 21341 2451
rect 21343 2445 21415 2451
rect 21525 2451 21815 2479
rect 21925 2469 22217 2497
rect 22349 2479 22375 2513
rect 21925 2463 21941 2469
rect 21525 2445 21541 2451
rect 19983 2128 20017 2420
rect 20141 2411 20415 2420
rect 20543 2411 20575 2445
rect 20583 2411 20615 2445
rect 20743 2411 20775 2445
rect 20783 2411 20815 2445
rect 20943 2411 20975 2445
rect 20983 2411 21015 2445
rect 21143 2411 21175 2445
rect 21183 2411 21215 2445
rect 21343 2411 21375 2445
rect 21383 2411 21415 2445
rect 21543 2420 21815 2451
rect 21943 2461 22217 2469
rect 21943 2420 22215 2461
rect 22325 2451 22375 2479
rect 22383 2461 22417 2513
rect 22549 2479 22575 2513
rect 22383 2451 22415 2461
rect 22325 2445 22341 2451
rect 22343 2445 22415 2451
rect 22525 2451 22575 2479
rect 22583 2461 22617 2513
rect 22749 2479 22775 2513
rect 22583 2451 22615 2461
rect 22525 2445 22541 2451
rect 22543 2445 22615 2451
rect 22725 2451 22775 2479
rect 22783 2461 22817 2513
rect 22949 2479 22975 2513
rect 22783 2451 22815 2461
rect 22725 2445 22741 2451
rect 22743 2445 22815 2451
rect 22925 2451 22975 2479
rect 22983 2461 23017 2513
rect 23149 2479 23175 2513
rect 22983 2451 23015 2461
rect 22925 2445 22941 2451
rect 22943 2445 23015 2451
rect 23125 2451 23175 2479
rect 23183 2461 23217 2513
rect 23347 2479 23617 2513
rect 23747 2513 25417 2531
rect 23747 2497 24017 2513
rect 23183 2451 23215 2461
rect 23125 2445 23141 2451
rect 23143 2445 23215 2451
rect 23325 2451 23615 2479
rect 23725 2469 24017 2497
rect 24149 2479 24175 2513
rect 23725 2463 23741 2469
rect 23325 2445 23341 2451
rect 21543 2411 21817 2420
rect 20027 2162 20051 2386
rect 20107 2382 20131 2386
rect 20059 2178 20061 2370
rect 20063 2166 20067 2382
rect 20085 2166 20131 2382
rect 20107 2162 20131 2166
rect 20141 2153 20417 2411
rect 20541 2405 20617 2411
rect 20427 2153 20451 2377
rect 20507 2373 20531 2377
rect 20459 2169 20461 2361
rect 20463 2157 20467 2373
rect 20485 2157 20531 2373
rect 20507 2153 20531 2157
rect 20541 2153 20575 2405
rect 20125 2128 20417 2153
rect 19983 2125 20015 2128
rect 19943 2119 20015 2125
rect 20125 2119 20141 2128
rect 20143 2119 20417 2128
rect 20525 2125 20575 2153
rect 20583 2125 20617 2405
rect 20741 2405 20817 2411
rect 20627 2153 20651 2377
rect 20707 2373 20731 2377
rect 20659 2169 20661 2361
rect 20663 2157 20667 2373
rect 20685 2157 20731 2373
rect 20707 2153 20731 2157
rect 20741 2153 20775 2405
rect 20525 2119 20617 2125
rect 20725 2125 20775 2153
rect 20783 2125 20817 2405
rect 20941 2405 21017 2411
rect 20827 2153 20851 2377
rect 20907 2373 20931 2377
rect 20859 2169 20861 2361
rect 20863 2157 20867 2373
rect 20885 2157 20931 2373
rect 20907 2153 20931 2157
rect 20941 2153 20975 2405
rect 20725 2119 20817 2125
rect 20925 2125 20975 2153
rect 20983 2125 21017 2405
rect 21141 2405 21217 2411
rect 21027 2153 21051 2377
rect 21107 2373 21131 2377
rect 21059 2169 21061 2361
rect 21063 2157 21067 2373
rect 21085 2157 21131 2373
rect 21107 2153 21131 2157
rect 21141 2153 21175 2405
rect 20925 2119 21017 2125
rect 21125 2125 21175 2153
rect 21183 2125 21217 2405
rect 21341 2405 21417 2411
rect 21227 2153 21251 2377
rect 21307 2373 21331 2377
rect 21259 2169 21261 2361
rect 21263 2157 21267 2373
rect 21285 2157 21331 2373
rect 21307 2153 21331 2157
rect 21341 2153 21375 2405
rect 21125 2119 21217 2125
rect 21325 2125 21375 2153
rect 21383 2125 21417 2405
rect 21427 2153 21451 2377
rect 21507 2373 21531 2377
rect 21459 2169 21461 2361
rect 21463 2157 21467 2373
rect 21485 2157 21531 2373
rect 21507 2153 21531 2157
rect 21541 2153 21817 2411
rect 21941 2411 22215 2420
rect 22343 2411 22375 2445
rect 22383 2411 22415 2445
rect 22543 2411 22575 2445
rect 22583 2411 22615 2445
rect 22743 2411 22775 2445
rect 22783 2411 22815 2445
rect 22943 2411 22975 2445
rect 22983 2411 23015 2445
rect 23143 2411 23175 2445
rect 23183 2411 23215 2445
rect 23343 2420 23615 2451
rect 23743 2461 24017 2469
rect 23743 2420 24015 2461
rect 24125 2451 24175 2479
rect 24183 2461 24217 2513
rect 24349 2479 24375 2513
rect 24183 2451 24215 2461
rect 24125 2445 24141 2451
rect 24143 2445 24215 2451
rect 24325 2451 24375 2479
rect 24383 2461 24417 2513
rect 24549 2479 24575 2513
rect 24383 2451 24415 2461
rect 24325 2445 24341 2451
rect 24343 2445 24415 2451
rect 24525 2451 24575 2479
rect 24583 2461 24617 2513
rect 24749 2479 24775 2513
rect 24583 2451 24615 2461
rect 24525 2445 24541 2451
rect 24543 2445 24615 2451
rect 24725 2451 24775 2479
rect 24783 2461 24817 2513
rect 24949 2479 24975 2513
rect 24783 2451 24815 2461
rect 24725 2445 24741 2451
rect 24743 2445 24815 2451
rect 24925 2451 24975 2479
rect 24983 2461 25017 2513
rect 25147 2479 25417 2513
rect 25547 2513 27217 2531
rect 25547 2497 25817 2513
rect 24983 2451 25015 2461
rect 24925 2445 24941 2451
rect 24943 2445 25015 2451
rect 25125 2451 25415 2479
rect 25525 2469 25817 2497
rect 25949 2479 25975 2513
rect 25525 2463 25541 2469
rect 25125 2445 25141 2451
rect 23343 2411 23617 2420
rect 21827 2162 21851 2386
rect 21907 2382 21931 2386
rect 21859 2178 21861 2370
rect 21863 2166 21867 2382
rect 21885 2166 21931 2382
rect 21907 2162 21931 2166
rect 21941 2153 22217 2411
rect 22341 2405 22417 2411
rect 22227 2153 22251 2377
rect 22307 2373 22331 2377
rect 22259 2169 22261 2361
rect 22263 2157 22267 2373
rect 22285 2157 22331 2373
rect 22307 2153 22331 2157
rect 22341 2153 22375 2405
rect 21325 2119 21417 2125
rect 21525 2128 21817 2153
rect 21925 2128 22217 2153
rect 21525 2119 21815 2128
rect 21925 2119 21941 2128
rect 21943 2119 22217 2128
rect 22325 2125 22375 2153
rect 22383 2125 22417 2405
rect 22541 2405 22617 2411
rect 22427 2153 22451 2377
rect 22507 2373 22531 2377
rect 22459 2169 22461 2361
rect 22463 2157 22467 2373
rect 22485 2157 22531 2373
rect 22507 2153 22531 2157
rect 22541 2153 22575 2405
rect 22325 2119 22417 2125
rect 22525 2125 22575 2153
rect 22583 2125 22617 2405
rect 22741 2405 22817 2411
rect 22627 2153 22651 2377
rect 22707 2373 22731 2377
rect 22659 2169 22661 2361
rect 22663 2157 22667 2373
rect 22685 2157 22731 2373
rect 22707 2153 22731 2157
rect 22741 2153 22775 2405
rect 22525 2119 22617 2125
rect 22725 2125 22775 2153
rect 22783 2125 22817 2405
rect 22941 2405 23017 2411
rect 22827 2153 22851 2377
rect 22907 2373 22931 2377
rect 22859 2169 22861 2361
rect 22863 2157 22867 2373
rect 22885 2157 22931 2373
rect 22907 2153 22931 2157
rect 22941 2153 22975 2405
rect 22725 2119 22817 2125
rect 22925 2125 22975 2153
rect 22983 2125 23017 2405
rect 23141 2405 23217 2411
rect 23027 2153 23051 2377
rect 23107 2373 23131 2377
rect 23059 2169 23061 2361
rect 23063 2157 23067 2373
rect 23085 2157 23131 2373
rect 23107 2153 23131 2157
rect 23141 2153 23175 2405
rect 22925 2119 23017 2125
rect 23125 2125 23175 2153
rect 23183 2125 23217 2405
rect 23227 2153 23251 2377
rect 23307 2373 23331 2377
rect 23259 2169 23261 2361
rect 23263 2157 23267 2373
rect 23285 2157 23331 2373
rect 23307 2153 23331 2157
rect 23341 2153 23617 2411
rect 23741 2411 24015 2420
rect 24143 2411 24175 2445
rect 24183 2411 24215 2445
rect 24343 2411 24375 2445
rect 24383 2411 24415 2445
rect 24543 2411 24575 2445
rect 24583 2411 24615 2445
rect 24743 2411 24775 2445
rect 24783 2411 24815 2445
rect 24943 2411 24975 2445
rect 24983 2411 25015 2445
rect 25143 2420 25415 2451
rect 25543 2461 25817 2469
rect 25543 2420 25815 2461
rect 25925 2451 25975 2479
rect 25983 2461 26017 2513
rect 26149 2479 26175 2513
rect 25983 2451 26015 2461
rect 25925 2445 25941 2451
rect 25943 2445 26015 2451
rect 26125 2451 26175 2479
rect 26183 2461 26217 2513
rect 26349 2479 26375 2513
rect 26183 2451 26215 2461
rect 26125 2445 26141 2451
rect 26143 2445 26215 2451
rect 26325 2451 26375 2479
rect 26383 2461 26417 2513
rect 26549 2479 26575 2513
rect 26383 2451 26415 2461
rect 26325 2445 26341 2451
rect 26343 2445 26415 2451
rect 26525 2451 26575 2479
rect 26583 2461 26617 2513
rect 26749 2479 26775 2513
rect 26583 2451 26615 2461
rect 26525 2445 26541 2451
rect 26543 2445 26615 2451
rect 26725 2451 26775 2479
rect 26783 2461 26817 2513
rect 26947 2479 27217 2513
rect 27347 2513 29017 2531
rect 27347 2497 27617 2513
rect 26783 2451 26815 2461
rect 26725 2445 26741 2451
rect 26743 2445 26815 2451
rect 26925 2451 27215 2479
rect 27325 2469 27617 2497
rect 27749 2479 27775 2513
rect 27325 2463 27341 2469
rect 26925 2445 26941 2451
rect 25143 2411 25417 2420
rect 23627 2162 23651 2386
rect 23707 2382 23731 2386
rect 23659 2178 23661 2370
rect 23663 2166 23667 2382
rect 23685 2166 23731 2382
rect 23707 2162 23731 2166
rect 23741 2153 24017 2411
rect 24141 2405 24217 2411
rect 24027 2153 24051 2377
rect 24107 2373 24131 2377
rect 24059 2169 24061 2361
rect 24063 2157 24067 2373
rect 24085 2157 24131 2373
rect 24107 2153 24131 2157
rect 24141 2153 24175 2405
rect 23125 2119 23217 2125
rect 23325 2128 23617 2153
rect 23725 2128 24017 2153
rect 23325 2119 23615 2128
rect 23725 2119 23741 2128
rect 23743 2119 24017 2128
rect 24125 2125 24175 2153
rect 24183 2125 24217 2405
rect 24341 2405 24417 2411
rect 24227 2153 24251 2377
rect 24307 2373 24331 2377
rect 24259 2169 24261 2361
rect 24263 2157 24267 2373
rect 24285 2157 24331 2373
rect 24307 2153 24331 2157
rect 24341 2153 24375 2405
rect 24125 2119 24217 2125
rect 24325 2125 24375 2153
rect 24383 2125 24417 2405
rect 24541 2405 24617 2411
rect 24427 2153 24451 2377
rect 24507 2373 24531 2377
rect 24459 2169 24461 2361
rect 24463 2157 24467 2373
rect 24485 2157 24531 2373
rect 24507 2153 24531 2157
rect 24541 2153 24575 2405
rect 24325 2119 24417 2125
rect 24525 2125 24575 2153
rect 24583 2125 24617 2405
rect 24741 2405 24817 2411
rect 24627 2153 24651 2377
rect 24707 2373 24731 2377
rect 24659 2169 24661 2361
rect 24663 2157 24667 2373
rect 24685 2157 24731 2373
rect 24707 2153 24731 2157
rect 24741 2153 24775 2405
rect 24525 2119 24617 2125
rect 24725 2125 24775 2153
rect 24783 2125 24817 2405
rect 24941 2405 25017 2411
rect 24827 2153 24851 2377
rect 24907 2373 24931 2377
rect 24859 2169 24861 2361
rect 24863 2157 24867 2373
rect 24885 2157 24931 2373
rect 24907 2153 24931 2157
rect 24941 2153 24975 2405
rect 24725 2119 24817 2125
rect 24925 2125 24975 2153
rect 24983 2125 25017 2405
rect 25027 2153 25051 2377
rect 25107 2373 25131 2377
rect 25059 2169 25061 2361
rect 25063 2157 25067 2373
rect 25085 2157 25131 2373
rect 25107 2153 25131 2157
rect 25141 2153 25417 2411
rect 25541 2411 25815 2420
rect 25943 2411 25975 2445
rect 25983 2411 26015 2445
rect 26143 2411 26175 2445
rect 26183 2411 26215 2445
rect 26343 2411 26375 2445
rect 26383 2411 26415 2445
rect 26543 2411 26575 2445
rect 26583 2411 26615 2445
rect 26743 2411 26775 2445
rect 26783 2411 26815 2445
rect 26943 2420 27215 2451
rect 27343 2461 27617 2469
rect 27343 2420 27615 2461
rect 27725 2451 27775 2479
rect 27783 2461 27817 2513
rect 27949 2479 27975 2513
rect 27783 2451 27815 2461
rect 27725 2445 27741 2451
rect 27743 2445 27815 2451
rect 27925 2451 27975 2479
rect 27983 2461 28017 2513
rect 28149 2479 28175 2513
rect 27983 2451 28015 2461
rect 27925 2445 27941 2451
rect 27943 2445 28015 2451
rect 28125 2451 28175 2479
rect 28183 2461 28217 2513
rect 28349 2479 28375 2513
rect 28183 2451 28215 2461
rect 28125 2445 28141 2451
rect 28143 2445 28215 2451
rect 28325 2451 28375 2479
rect 28383 2461 28417 2513
rect 28549 2479 28575 2513
rect 28383 2451 28415 2461
rect 28325 2445 28341 2451
rect 28343 2445 28415 2451
rect 28525 2451 28575 2479
rect 28583 2461 28617 2513
rect 28747 2479 29017 2513
rect 29147 2513 30817 2531
rect 29147 2497 29417 2513
rect 28583 2451 28615 2461
rect 28525 2445 28541 2451
rect 28543 2445 28615 2451
rect 28725 2451 29015 2479
rect 29125 2469 29417 2497
rect 29549 2479 29575 2513
rect 29125 2463 29141 2469
rect 28725 2445 28741 2451
rect 26943 2411 27217 2420
rect 25427 2162 25451 2386
rect 25507 2382 25531 2386
rect 25459 2178 25461 2370
rect 25463 2166 25467 2382
rect 25485 2166 25531 2382
rect 25507 2162 25531 2166
rect 25541 2153 25817 2411
rect 25941 2405 26017 2411
rect 25827 2153 25851 2377
rect 25907 2373 25931 2377
rect 25859 2169 25861 2361
rect 25863 2157 25867 2373
rect 25885 2157 25931 2373
rect 25907 2153 25931 2157
rect 25941 2153 25975 2405
rect 24925 2119 25017 2125
rect 25125 2128 25417 2153
rect 25525 2128 25817 2153
rect 25125 2119 25415 2128
rect 25525 2119 25541 2128
rect 25543 2119 25817 2128
rect 25925 2125 25975 2153
rect 25983 2125 26017 2405
rect 26141 2405 26217 2411
rect 26027 2153 26051 2377
rect 26107 2373 26131 2377
rect 26059 2169 26061 2361
rect 26063 2157 26067 2373
rect 26085 2157 26131 2373
rect 26107 2153 26131 2157
rect 26141 2153 26175 2405
rect 25925 2119 26017 2125
rect 26125 2125 26175 2153
rect 26183 2125 26217 2405
rect 26341 2405 26417 2411
rect 26227 2153 26251 2377
rect 26307 2373 26331 2377
rect 26259 2169 26261 2361
rect 26263 2157 26267 2373
rect 26285 2157 26331 2373
rect 26307 2153 26331 2157
rect 26341 2153 26375 2405
rect 26125 2119 26217 2125
rect 26325 2125 26375 2153
rect 26383 2125 26417 2405
rect 26541 2405 26617 2411
rect 26427 2153 26451 2377
rect 26507 2373 26531 2377
rect 26459 2169 26461 2361
rect 26463 2157 26467 2373
rect 26485 2157 26531 2373
rect 26507 2153 26531 2157
rect 26541 2153 26575 2405
rect 26325 2119 26417 2125
rect 26525 2125 26575 2153
rect 26583 2125 26617 2405
rect 26741 2405 26817 2411
rect 26627 2153 26651 2377
rect 26707 2373 26731 2377
rect 26659 2169 26661 2361
rect 26663 2157 26667 2373
rect 26685 2157 26731 2373
rect 26707 2153 26731 2157
rect 26741 2153 26775 2405
rect 26525 2119 26617 2125
rect 26725 2125 26775 2153
rect 26783 2125 26817 2405
rect 26827 2153 26851 2377
rect 26907 2373 26931 2377
rect 26859 2169 26861 2361
rect 26863 2157 26867 2373
rect 26885 2157 26931 2373
rect 26907 2153 26931 2157
rect 26941 2153 27217 2411
rect 27341 2411 27615 2420
rect 27743 2411 27775 2445
rect 27783 2411 27815 2445
rect 27943 2411 27975 2445
rect 27983 2411 28015 2445
rect 28143 2411 28175 2445
rect 28183 2411 28215 2445
rect 28343 2411 28375 2445
rect 28383 2411 28415 2445
rect 28543 2411 28575 2445
rect 28583 2411 28615 2445
rect 28743 2420 29015 2451
rect 29143 2461 29417 2469
rect 29143 2420 29415 2461
rect 29525 2451 29575 2479
rect 29583 2461 29617 2513
rect 29749 2479 29775 2513
rect 29583 2451 29615 2461
rect 29525 2445 29541 2451
rect 29543 2445 29615 2451
rect 29725 2451 29775 2479
rect 29783 2461 29817 2513
rect 29949 2479 29975 2513
rect 29783 2451 29815 2461
rect 29725 2445 29741 2451
rect 29743 2445 29815 2451
rect 29925 2451 29975 2479
rect 29983 2461 30017 2513
rect 30149 2479 30175 2513
rect 29983 2451 30015 2461
rect 29925 2445 29941 2451
rect 29943 2445 30015 2451
rect 30125 2451 30175 2479
rect 30183 2461 30217 2513
rect 30349 2479 30375 2513
rect 30183 2451 30215 2461
rect 30125 2445 30141 2451
rect 30143 2445 30215 2451
rect 30325 2451 30375 2479
rect 30383 2461 30417 2513
rect 30547 2479 30817 2513
rect 30947 2513 32617 2531
rect 30947 2497 31217 2513
rect 30383 2451 30415 2461
rect 30325 2445 30341 2451
rect 30343 2445 30415 2451
rect 30525 2451 30815 2479
rect 30925 2469 31217 2497
rect 31349 2479 31375 2513
rect 30925 2463 30941 2469
rect 30525 2445 30541 2451
rect 28743 2411 29017 2420
rect 27227 2162 27251 2386
rect 27307 2382 27331 2386
rect 27259 2178 27261 2370
rect 27263 2166 27267 2382
rect 27285 2166 27331 2382
rect 27307 2162 27331 2166
rect 27341 2153 27617 2411
rect 27741 2405 27817 2411
rect 27627 2153 27651 2377
rect 27707 2373 27731 2377
rect 27659 2169 27661 2361
rect 27663 2157 27667 2373
rect 27685 2157 27731 2373
rect 27707 2153 27731 2157
rect 27741 2153 27775 2405
rect 26725 2119 26817 2125
rect 26925 2128 27217 2153
rect 27325 2128 27617 2153
rect 26925 2119 27215 2128
rect 27325 2119 27341 2128
rect 27343 2119 27617 2128
rect 27725 2125 27775 2153
rect 27783 2125 27817 2405
rect 27941 2405 28017 2411
rect 27827 2153 27851 2377
rect 27907 2373 27931 2377
rect 27859 2169 27861 2361
rect 27863 2157 27867 2373
rect 27885 2157 27931 2373
rect 27907 2153 27931 2157
rect 27941 2153 27975 2405
rect 27725 2119 27817 2125
rect 27925 2125 27975 2153
rect 27983 2125 28017 2405
rect 28141 2405 28217 2411
rect 28027 2153 28051 2377
rect 28107 2373 28131 2377
rect 28059 2169 28061 2361
rect 28063 2157 28067 2373
rect 28085 2157 28131 2373
rect 28107 2153 28131 2157
rect 28141 2153 28175 2405
rect 27925 2119 28017 2125
rect 28125 2125 28175 2153
rect 28183 2125 28217 2405
rect 28341 2405 28417 2411
rect 28227 2153 28251 2377
rect 28307 2373 28331 2377
rect 28259 2169 28261 2361
rect 28263 2157 28267 2373
rect 28285 2157 28331 2373
rect 28307 2153 28331 2157
rect 28341 2153 28375 2405
rect 28125 2119 28217 2125
rect 28325 2125 28375 2153
rect 28383 2125 28417 2405
rect 28541 2405 28617 2411
rect 28427 2153 28451 2377
rect 28507 2373 28531 2377
rect 28459 2169 28461 2361
rect 28463 2157 28467 2373
rect 28485 2157 28531 2373
rect 28507 2153 28531 2157
rect 28541 2153 28575 2405
rect 28325 2119 28417 2125
rect 28525 2125 28575 2153
rect 28583 2125 28617 2405
rect 28627 2153 28651 2377
rect 28707 2373 28731 2377
rect 28659 2169 28661 2361
rect 28663 2157 28667 2373
rect 28685 2157 28731 2373
rect 28707 2153 28731 2157
rect 28741 2153 29017 2411
rect 29141 2411 29415 2420
rect 29543 2411 29575 2445
rect 29583 2411 29615 2445
rect 29743 2411 29775 2445
rect 29783 2411 29815 2445
rect 29943 2411 29975 2445
rect 29983 2411 30015 2445
rect 30143 2411 30175 2445
rect 30183 2411 30215 2445
rect 30343 2411 30375 2445
rect 30383 2411 30415 2445
rect 30543 2420 30815 2451
rect 30943 2461 31217 2469
rect 30943 2420 31215 2461
rect 31325 2451 31375 2479
rect 31383 2461 31417 2513
rect 31549 2479 31575 2513
rect 31383 2451 31415 2461
rect 31325 2445 31341 2451
rect 31343 2445 31415 2451
rect 31525 2451 31575 2479
rect 31583 2461 31617 2513
rect 31749 2479 31775 2513
rect 31583 2451 31615 2461
rect 31525 2445 31541 2451
rect 31543 2445 31615 2451
rect 31725 2451 31775 2479
rect 31783 2461 31817 2513
rect 31949 2479 31975 2513
rect 31783 2451 31815 2461
rect 31725 2445 31741 2451
rect 31743 2445 31815 2451
rect 31925 2451 31975 2479
rect 31983 2461 32017 2513
rect 32149 2479 32175 2513
rect 31983 2451 32015 2461
rect 31925 2445 31941 2451
rect 31943 2445 32015 2451
rect 32125 2451 32175 2479
rect 32183 2461 32217 2513
rect 32347 2479 32617 2513
rect 32747 2513 34417 2531
rect 32747 2497 33017 2513
rect 32183 2451 32215 2461
rect 32125 2445 32141 2451
rect 32143 2445 32215 2451
rect 32325 2451 32615 2479
rect 32725 2469 33017 2497
rect 33149 2479 33175 2513
rect 32725 2463 32741 2469
rect 32325 2445 32341 2451
rect 30543 2411 30817 2420
rect 29027 2162 29051 2386
rect 29107 2382 29131 2386
rect 29059 2178 29061 2370
rect 29063 2166 29067 2382
rect 29085 2166 29131 2382
rect 29107 2162 29131 2166
rect 29141 2153 29417 2411
rect 29541 2405 29617 2411
rect 29427 2153 29451 2377
rect 29507 2373 29531 2377
rect 29459 2169 29461 2361
rect 29463 2157 29467 2373
rect 29485 2157 29531 2373
rect 29507 2153 29531 2157
rect 29541 2153 29575 2405
rect 28525 2119 28617 2125
rect 28725 2128 29017 2153
rect 29125 2128 29417 2153
rect 28725 2119 29015 2128
rect 29125 2119 29141 2128
rect 29143 2119 29417 2128
rect 29525 2125 29575 2153
rect 29583 2125 29617 2405
rect 29741 2405 29817 2411
rect 29627 2153 29651 2377
rect 29707 2373 29731 2377
rect 29659 2169 29661 2361
rect 29663 2157 29667 2373
rect 29685 2157 29731 2373
rect 29707 2153 29731 2157
rect 29741 2153 29775 2405
rect 29525 2119 29617 2125
rect 29725 2125 29775 2153
rect 29783 2125 29817 2405
rect 29941 2405 30017 2411
rect 29827 2153 29851 2377
rect 29907 2373 29931 2377
rect 29859 2169 29861 2361
rect 29863 2157 29867 2373
rect 29885 2157 29931 2373
rect 29907 2153 29931 2157
rect 29941 2153 29975 2405
rect 29725 2119 29817 2125
rect 29925 2125 29975 2153
rect 29983 2125 30017 2405
rect 30141 2405 30217 2411
rect 30027 2153 30051 2377
rect 30107 2373 30131 2377
rect 30059 2169 30061 2361
rect 30063 2157 30067 2373
rect 30085 2157 30131 2373
rect 30107 2153 30131 2157
rect 30141 2153 30175 2405
rect 29925 2119 30017 2125
rect 30125 2125 30175 2153
rect 30183 2125 30217 2405
rect 30341 2405 30417 2411
rect 30227 2153 30251 2377
rect 30307 2373 30331 2377
rect 30259 2169 30261 2361
rect 30263 2157 30267 2373
rect 30285 2157 30331 2373
rect 30307 2153 30331 2157
rect 30341 2153 30375 2405
rect 30125 2119 30217 2125
rect 30325 2125 30375 2153
rect 30383 2125 30417 2405
rect 30427 2153 30451 2377
rect 30507 2373 30531 2377
rect 30459 2169 30461 2361
rect 30463 2157 30467 2373
rect 30485 2157 30531 2373
rect 30507 2153 30531 2157
rect 30541 2153 30817 2411
rect 30941 2411 31215 2420
rect 31343 2411 31375 2445
rect 31383 2411 31415 2445
rect 31543 2411 31575 2445
rect 31583 2411 31615 2445
rect 31743 2411 31775 2445
rect 31783 2411 31815 2445
rect 31943 2411 31975 2445
rect 31983 2411 32015 2445
rect 32143 2411 32175 2445
rect 32183 2411 32215 2445
rect 32343 2420 32615 2451
rect 32743 2461 33017 2469
rect 32743 2420 33015 2461
rect 33125 2451 33175 2479
rect 33183 2461 33217 2513
rect 33349 2479 33375 2513
rect 33183 2451 33215 2461
rect 33125 2445 33141 2451
rect 33143 2445 33215 2451
rect 33325 2451 33375 2479
rect 33383 2461 33417 2513
rect 33549 2479 33575 2513
rect 33383 2451 33415 2461
rect 33325 2445 33341 2451
rect 33343 2445 33415 2451
rect 33525 2451 33575 2479
rect 33583 2461 33617 2513
rect 33749 2479 33775 2513
rect 33583 2451 33615 2461
rect 33525 2445 33541 2451
rect 33543 2445 33615 2451
rect 33725 2451 33775 2479
rect 33783 2461 33817 2513
rect 33949 2479 33975 2513
rect 33783 2451 33815 2461
rect 33725 2445 33741 2451
rect 33743 2445 33815 2451
rect 33925 2451 33975 2479
rect 33983 2461 34017 2513
rect 34147 2479 34417 2513
rect 34547 2513 36217 2531
rect 34547 2497 34817 2513
rect 33983 2451 34015 2461
rect 33925 2445 33941 2451
rect 33943 2445 34015 2451
rect 34125 2451 34415 2479
rect 34525 2469 34817 2497
rect 34949 2479 34975 2513
rect 34525 2463 34541 2469
rect 34125 2445 34141 2451
rect 32343 2411 32617 2420
rect 30827 2162 30851 2386
rect 30907 2382 30931 2386
rect 30859 2178 30861 2370
rect 30863 2166 30867 2382
rect 30885 2166 30931 2382
rect 30907 2162 30931 2166
rect 30941 2153 31217 2411
rect 31341 2405 31417 2411
rect 31227 2153 31251 2377
rect 31307 2373 31331 2377
rect 31259 2169 31261 2361
rect 31263 2157 31267 2373
rect 31285 2157 31331 2373
rect 31307 2153 31331 2157
rect 31341 2153 31375 2405
rect 30325 2119 30417 2125
rect 30525 2128 30817 2153
rect 30925 2128 31217 2153
rect 30525 2119 30815 2128
rect 30925 2119 30941 2128
rect 30943 2119 31217 2128
rect 31325 2125 31375 2153
rect 31383 2125 31417 2405
rect 31541 2405 31617 2411
rect 31427 2153 31451 2377
rect 31507 2373 31531 2377
rect 31459 2169 31461 2361
rect 31463 2157 31467 2373
rect 31485 2157 31531 2373
rect 31507 2153 31531 2157
rect 31541 2153 31575 2405
rect 31325 2119 31417 2125
rect 31525 2125 31575 2153
rect 31583 2125 31617 2405
rect 31741 2405 31817 2411
rect 31627 2153 31651 2377
rect 31707 2373 31731 2377
rect 31659 2169 31661 2361
rect 31663 2157 31667 2373
rect 31685 2157 31731 2373
rect 31707 2153 31731 2157
rect 31741 2153 31775 2405
rect 31525 2119 31617 2125
rect 31725 2125 31775 2153
rect 31783 2125 31817 2405
rect 31941 2405 32017 2411
rect 31827 2153 31851 2377
rect 31907 2373 31931 2377
rect 31859 2169 31861 2361
rect 31863 2157 31867 2373
rect 31885 2157 31931 2373
rect 31907 2153 31931 2157
rect 31941 2153 31975 2405
rect 31725 2119 31817 2125
rect 31925 2125 31975 2153
rect 31983 2125 32017 2405
rect 32141 2405 32217 2411
rect 32027 2153 32051 2377
rect 32107 2373 32131 2377
rect 32059 2169 32061 2361
rect 32063 2157 32067 2373
rect 32085 2157 32131 2373
rect 32107 2153 32131 2157
rect 32141 2153 32175 2405
rect 31925 2119 32017 2125
rect 32125 2125 32175 2153
rect 32183 2125 32217 2405
rect 32227 2153 32251 2377
rect 32307 2373 32331 2377
rect 32259 2169 32261 2361
rect 32263 2157 32267 2373
rect 32285 2157 32331 2373
rect 32307 2153 32331 2157
rect 32341 2153 32617 2411
rect 32741 2411 33015 2420
rect 33143 2411 33175 2445
rect 33183 2411 33215 2445
rect 33343 2411 33375 2445
rect 33383 2411 33415 2445
rect 33543 2411 33575 2445
rect 33583 2411 33615 2445
rect 33743 2411 33775 2445
rect 33783 2411 33815 2445
rect 33943 2411 33975 2445
rect 33983 2411 34015 2445
rect 34143 2420 34415 2451
rect 34543 2461 34817 2469
rect 34543 2420 34815 2461
rect 34925 2451 34975 2479
rect 34983 2461 35017 2513
rect 35149 2479 35175 2513
rect 34983 2451 35015 2461
rect 34925 2445 34941 2451
rect 34943 2445 35015 2451
rect 35125 2451 35175 2479
rect 35183 2461 35217 2513
rect 35349 2479 35375 2513
rect 35183 2451 35215 2461
rect 35125 2445 35141 2451
rect 35143 2445 35215 2451
rect 35325 2451 35375 2479
rect 35383 2461 35417 2513
rect 35549 2479 35575 2513
rect 35383 2451 35415 2461
rect 35325 2445 35341 2451
rect 35343 2445 35415 2451
rect 35525 2451 35575 2479
rect 35583 2461 35617 2513
rect 35749 2479 35775 2513
rect 35583 2451 35615 2461
rect 35525 2445 35541 2451
rect 35543 2445 35615 2451
rect 35725 2451 35775 2479
rect 35783 2461 35817 2513
rect 35947 2479 36217 2513
rect 36347 2513 38017 2531
rect 36347 2497 36617 2513
rect 35783 2451 35815 2461
rect 35725 2445 35741 2451
rect 35743 2445 35815 2451
rect 35925 2451 36215 2479
rect 36325 2469 36617 2497
rect 36749 2479 36775 2513
rect 36325 2463 36341 2469
rect 35925 2445 35941 2451
rect 34143 2411 34417 2420
rect 32627 2162 32651 2386
rect 32707 2382 32731 2386
rect 32659 2178 32661 2370
rect 32663 2166 32667 2382
rect 32685 2166 32731 2382
rect 32707 2162 32731 2166
rect 32741 2153 33017 2411
rect 33141 2405 33217 2411
rect 33027 2153 33051 2377
rect 33107 2373 33131 2377
rect 33059 2169 33061 2361
rect 33063 2157 33067 2373
rect 33085 2157 33131 2373
rect 33107 2153 33131 2157
rect 33141 2153 33175 2405
rect 32125 2119 32217 2125
rect 32325 2128 32617 2153
rect 32725 2128 33017 2153
rect 32325 2119 32615 2128
rect 32725 2119 32741 2128
rect 32743 2119 33017 2128
rect 33125 2125 33175 2153
rect 33183 2125 33217 2405
rect 33341 2405 33417 2411
rect 33227 2153 33251 2377
rect 33307 2373 33331 2377
rect 33259 2169 33261 2361
rect 33263 2157 33267 2373
rect 33285 2157 33331 2373
rect 33307 2153 33331 2157
rect 33341 2153 33375 2405
rect 33125 2119 33217 2125
rect 33325 2125 33375 2153
rect 33383 2125 33417 2405
rect 33541 2405 33617 2411
rect 33427 2153 33451 2377
rect 33507 2373 33531 2377
rect 33459 2169 33461 2361
rect 33463 2157 33467 2373
rect 33485 2157 33531 2373
rect 33507 2153 33531 2157
rect 33541 2153 33575 2405
rect 33325 2119 33417 2125
rect 33525 2125 33575 2153
rect 33583 2125 33617 2405
rect 33741 2405 33817 2411
rect 33627 2153 33651 2377
rect 33707 2373 33731 2377
rect 33659 2169 33661 2361
rect 33663 2157 33667 2373
rect 33685 2157 33731 2373
rect 33707 2153 33731 2157
rect 33741 2153 33775 2405
rect 33525 2119 33617 2125
rect 33725 2125 33775 2153
rect 33783 2125 33817 2405
rect 33941 2405 34017 2411
rect 33827 2153 33851 2377
rect 33907 2373 33931 2377
rect 33859 2169 33861 2361
rect 33863 2157 33867 2373
rect 33885 2157 33931 2373
rect 33907 2153 33931 2157
rect 33941 2153 33975 2405
rect 33725 2119 33817 2125
rect 33925 2125 33975 2153
rect 33983 2125 34017 2405
rect 34027 2153 34051 2377
rect 34107 2373 34131 2377
rect 34059 2169 34061 2361
rect 34063 2157 34067 2373
rect 34085 2157 34131 2373
rect 34107 2153 34131 2157
rect 34141 2153 34417 2411
rect 34541 2411 34815 2420
rect 34943 2411 34975 2445
rect 34983 2411 35015 2445
rect 35143 2411 35175 2445
rect 35183 2411 35215 2445
rect 35343 2411 35375 2445
rect 35383 2411 35415 2445
rect 35543 2411 35575 2445
rect 35583 2411 35615 2445
rect 35743 2411 35775 2445
rect 35783 2411 35815 2445
rect 35943 2420 36215 2451
rect 36343 2461 36617 2469
rect 36343 2420 36615 2461
rect 36725 2451 36775 2479
rect 36783 2461 36817 2513
rect 36949 2479 36975 2513
rect 36783 2451 36815 2461
rect 36725 2445 36741 2451
rect 36743 2445 36815 2451
rect 36925 2451 36975 2479
rect 36983 2461 37017 2513
rect 37149 2479 37175 2513
rect 36983 2451 37015 2461
rect 36925 2445 36941 2451
rect 36943 2445 37015 2451
rect 37125 2451 37175 2479
rect 37183 2461 37217 2513
rect 37349 2479 37375 2513
rect 37183 2451 37215 2461
rect 37125 2445 37141 2451
rect 37143 2445 37215 2451
rect 37325 2451 37375 2479
rect 37383 2461 37417 2513
rect 37549 2479 37575 2513
rect 37383 2451 37415 2461
rect 37325 2445 37341 2451
rect 37343 2445 37415 2451
rect 37525 2451 37575 2479
rect 37583 2461 37617 2513
rect 37747 2479 38017 2513
rect 38147 2513 39817 2531
rect 38147 2497 38417 2513
rect 37583 2451 37615 2461
rect 37525 2445 37541 2451
rect 37543 2445 37615 2451
rect 37725 2451 38015 2479
rect 38125 2469 38417 2497
rect 38549 2479 38575 2513
rect 38125 2463 38141 2469
rect 37725 2445 37741 2451
rect 35943 2411 36217 2420
rect 34427 2162 34451 2386
rect 34507 2382 34531 2386
rect 34459 2178 34461 2370
rect 34463 2166 34467 2382
rect 34485 2166 34531 2382
rect 34507 2162 34531 2166
rect 34541 2153 34817 2411
rect 34941 2405 35017 2411
rect 34827 2153 34851 2377
rect 34907 2373 34931 2377
rect 34859 2169 34861 2361
rect 34863 2157 34867 2373
rect 34885 2157 34931 2373
rect 34907 2153 34931 2157
rect 34941 2153 34975 2405
rect 33925 2119 34017 2125
rect 34125 2128 34417 2153
rect 34525 2128 34817 2153
rect 34125 2119 34415 2128
rect 34525 2119 34541 2128
rect 34543 2119 34817 2128
rect 34925 2125 34975 2153
rect 34983 2125 35017 2405
rect 35141 2405 35217 2411
rect 35027 2153 35051 2377
rect 35107 2373 35131 2377
rect 35059 2169 35061 2361
rect 35063 2157 35067 2373
rect 35085 2157 35131 2373
rect 35107 2153 35131 2157
rect 35141 2153 35175 2405
rect 34925 2119 35017 2125
rect 35125 2125 35175 2153
rect 35183 2125 35217 2405
rect 35341 2405 35417 2411
rect 35227 2153 35251 2377
rect 35307 2373 35331 2377
rect 35259 2169 35261 2361
rect 35263 2157 35267 2373
rect 35285 2157 35331 2373
rect 35307 2153 35331 2157
rect 35341 2153 35375 2405
rect 35125 2119 35217 2125
rect 35325 2125 35375 2153
rect 35383 2125 35417 2405
rect 35541 2405 35617 2411
rect 35427 2153 35451 2377
rect 35507 2373 35531 2377
rect 35459 2169 35461 2361
rect 35463 2157 35467 2373
rect 35485 2157 35531 2373
rect 35507 2153 35531 2157
rect 35541 2153 35575 2405
rect 35325 2119 35417 2125
rect 35525 2125 35575 2153
rect 35583 2125 35617 2405
rect 35741 2405 35817 2411
rect 35627 2153 35651 2377
rect 35707 2373 35731 2377
rect 35659 2169 35661 2361
rect 35663 2157 35667 2373
rect 35685 2157 35731 2373
rect 35707 2153 35731 2157
rect 35741 2153 35775 2405
rect 35525 2119 35617 2125
rect 35725 2125 35775 2153
rect 35783 2125 35817 2405
rect 35827 2153 35851 2377
rect 35907 2373 35931 2377
rect 35859 2169 35861 2361
rect 35863 2157 35867 2373
rect 35885 2157 35931 2373
rect 35907 2153 35931 2157
rect 35941 2153 36217 2411
rect 36341 2411 36615 2420
rect 36743 2411 36775 2445
rect 36783 2411 36815 2445
rect 36943 2411 36975 2445
rect 36983 2411 37015 2445
rect 37143 2411 37175 2445
rect 37183 2411 37215 2445
rect 37343 2411 37375 2445
rect 37383 2411 37415 2445
rect 37543 2411 37575 2445
rect 37583 2411 37615 2445
rect 37743 2420 38015 2451
rect 38143 2461 38417 2469
rect 38143 2420 38415 2461
rect 38525 2451 38575 2479
rect 38583 2461 38617 2513
rect 38749 2479 38775 2513
rect 38583 2451 38615 2461
rect 38525 2445 38541 2451
rect 38543 2445 38615 2451
rect 38725 2451 38775 2479
rect 38783 2461 38817 2513
rect 38949 2479 38975 2513
rect 38783 2451 38815 2461
rect 38725 2445 38741 2451
rect 38743 2445 38815 2451
rect 38925 2451 38975 2479
rect 38983 2461 39017 2513
rect 39149 2479 39175 2513
rect 38983 2451 39015 2461
rect 38925 2445 38941 2451
rect 38943 2445 39015 2451
rect 39125 2451 39175 2479
rect 39183 2461 39217 2513
rect 39349 2479 39375 2513
rect 39183 2451 39215 2461
rect 39125 2445 39141 2451
rect 39143 2445 39215 2451
rect 39325 2451 39375 2479
rect 39383 2461 39417 2513
rect 39547 2479 39817 2513
rect 39947 2513 41617 2531
rect 39947 2497 40217 2513
rect 39383 2451 39415 2461
rect 39325 2445 39341 2451
rect 39343 2445 39415 2451
rect 39525 2451 39815 2479
rect 39925 2469 40217 2497
rect 40349 2479 40375 2513
rect 39925 2463 39941 2469
rect 39525 2445 39541 2451
rect 37743 2411 38017 2420
rect 36227 2162 36251 2386
rect 36307 2382 36331 2386
rect 36259 2178 36261 2370
rect 36263 2166 36267 2382
rect 36285 2166 36331 2382
rect 36307 2162 36331 2166
rect 36341 2153 36617 2411
rect 36741 2405 36817 2411
rect 36627 2153 36651 2377
rect 36707 2373 36731 2377
rect 36659 2169 36661 2361
rect 36663 2157 36667 2373
rect 36685 2157 36731 2373
rect 36707 2153 36731 2157
rect 36741 2153 36775 2405
rect 35725 2119 35817 2125
rect 35925 2128 36217 2153
rect 36325 2128 36617 2153
rect 35925 2119 36215 2128
rect 36325 2119 36341 2128
rect 36343 2119 36617 2128
rect 36725 2125 36775 2153
rect 36783 2125 36817 2405
rect 36941 2405 37017 2411
rect 36827 2153 36851 2377
rect 36907 2373 36931 2377
rect 36859 2169 36861 2361
rect 36863 2157 36867 2373
rect 36885 2157 36931 2373
rect 36907 2153 36931 2157
rect 36941 2153 36975 2405
rect 36725 2119 36817 2125
rect 36925 2125 36975 2153
rect 36983 2125 37017 2405
rect 37141 2405 37217 2411
rect 37027 2153 37051 2377
rect 37107 2373 37131 2377
rect 37059 2169 37061 2361
rect 37063 2157 37067 2373
rect 37085 2157 37131 2373
rect 37107 2153 37131 2157
rect 37141 2153 37175 2405
rect 36925 2119 37017 2125
rect 37125 2125 37175 2153
rect 37183 2125 37217 2405
rect 37341 2405 37417 2411
rect 37227 2153 37251 2377
rect 37307 2373 37331 2377
rect 37259 2169 37261 2361
rect 37263 2157 37267 2373
rect 37285 2157 37331 2373
rect 37307 2153 37331 2157
rect 37341 2153 37375 2405
rect 37125 2119 37217 2125
rect 37325 2125 37375 2153
rect 37383 2125 37417 2405
rect 37541 2405 37617 2411
rect 37427 2153 37451 2377
rect 37507 2373 37531 2377
rect 37459 2169 37461 2361
rect 37463 2157 37467 2373
rect 37485 2157 37531 2373
rect 37507 2153 37531 2157
rect 37541 2153 37575 2405
rect 37325 2119 37417 2125
rect 37525 2125 37575 2153
rect 37583 2125 37617 2405
rect 37627 2153 37651 2377
rect 37707 2373 37731 2377
rect 37659 2169 37661 2361
rect 37663 2157 37667 2373
rect 37685 2157 37731 2373
rect 37707 2153 37731 2157
rect 37741 2153 38017 2411
rect 38141 2411 38415 2420
rect 38543 2411 38575 2445
rect 38583 2411 38615 2445
rect 38743 2411 38775 2445
rect 38783 2411 38815 2445
rect 38943 2411 38975 2445
rect 38983 2411 39015 2445
rect 39143 2411 39175 2445
rect 39183 2411 39215 2445
rect 39343 2411 39375 2445
rect 39383 2411 39415 2445
rect 39543 2420 39815 2451
rect 39943 2461 40217 2469
rect 39943 2420 40215 2461
rect 40325 2451 40375 2479
rect 40383 2461 40417 2513
rect 40549 2479 40575 2513
rect 40383 2451 40415 2461
rect 40325 2445 40341 2451
rect 40343 2445 40415 2451
rect 40525 2451 40575 2479
rect 40583 2461 40617 2513
rect 40749 2479 40775 2513
rect 40583 2451 40615 2461
rect 40525 2445 40541 2451
rect 40543 2445 40615 2451
rect 40725 2451 40775 2479
rect 40783 2461 40817 2513
rect 40949 2479 40975 2513
rect 40783 2451 40815 2461
rect 40725 2445 40741 2451
rect 40743 2445 40815 2451
rect 40925 2451 40975 2479
rect 40983 2461 41017 2513
rect 41149 2479 41175 2513
rect 40983 2451 41015 2461
rect 40925 2445 40941 2451
rect 40943 2445 41015 2451
rect 41125 2451 41175 2479
rect 41183 2461 41217 2513
rect 41347 2479 41617 2513
rect 41747 2513 43417 2531
rect 41747 2497 42017 2513
rect 41183 2451 41215 2461
rect 41125 2445 41141 2451
rect 41143 2445 41215 2451
rect 41325 2451 41615 2479
rect 41725 2469 42017 2497
rect 42149 2479 42175 2513
rect 41725 2463 41741 2469
rect 41325 2445 41341 2451
rect 39543 2411 39817 2420
rect 38027 2162 38051 2386
rect 38107 2382 38131 2386
rect 38059 2178 38061 2370
rect 38063 2166 38067 2382
rect 38085 2166 38131 2382
rect 38107 2162 38131 2166
rect 38141 2153 38417 2411
rect 38541 2405 38617 2411
rect 38427 2153 38451 2377
rect 38507 2373 38531 2377
rect 38459 2169 38461 2361
rect 38463 2157 38467 2373
rect 38485 2157 38531 2373
rect 38507 2153 38531 2157
rect 38541 2153 38575 2405
rect 37525 2119 37617 2125
rect 37725 2128 38017 2153
rect 38125 2128 38417 2153
rect 37725 2119 38015 2128
rect 38125 2119 38141 2128
rect 38143 2119 38417 2128
rect 38525 2125 38575 2153
rect 38583 2125 38617 2405
rect 38741 2405 38817 2411
rect 38627 2153 38651 2377
rect 38707 2373 38731 2377
rect 38659 2169 38661 2361
rect 38663 2157 38667 2373
rect 38685 2157 38731 2373
rect 38707 2153 38731 2157
rect 38741 2153 38775 2405
rect 38525 2119 38617 2125
rect 38725 2125 38775 2153
rect 38783 2125 38817 2405
rect 38941 2405 39017 2411
rect 38827 2153 38851 2377
rect 38907 2373 38931 2377
rect 38859 2169 38861 2361
rect 38863 2157 38867 2373
rect 38885 2157 38931 2373
rect 38907 2153 38931 2157
rect 38941 2153 38975 2405
rect 38725 2119 38817 2125
rect 38925 2125 38975 2153
rect 38983 2125 39017 2405
rect 39141 2405 39217 2411
rect 39027 2153 39051 2377
rect 39107 2373 39131 2377
rect 39059 2169 39061 2361
rect 39063 2157 39067 2373
rect 39085 2157 39131 2373
rect 39107 2153 39131 2157
rect 39141 2153 39175 2405
rect 38925 2119 39017 2125
rect 39125 2125 39175 2153
rect 39183 2125 39217 2405
rect 39341 2405 39417 2411
rect 39227 2153 39251 2377
rect 39307 2373 39331 2377
rect 39259 2169 39261 2361
rect 39263 2157 39267 2373
rect 39285 2157 39331 2373
rect 39307 2153 39331 2157
rect 39341 2153 39375 2405
rect 39125 2119 39217 2125
rect 39325 2125 39375 2153
rect 39383 2125 39417 2405
rect 39427 2153 39451 2377
rect 39507 2373 39531 2377
rect 39459 2169 39461 2361
rect 39463 2157 39467 2373
rect 39485 2157 39531 2373
rect 39507 2153 39531 2157
rect 39541 2153 39817 2411
rect 39941 2411 40215 2420
rect 40343 2411 40375 2445
rect 40383 2411 40415 2445
rect 40543 2411 40575 2445
rect 40583 2411 40615 2445
rect 40743 2411 40775 2445
rect 40783 2411 40815 2445
rect 40943 2411 40975 2445
rect 40983 2411 41015 2445
rect 41143 2411 41175 2445
rect 41183 2411 41215 2445
rect 41343 2420 41615 2451
rect 41743 2461 42017 2469
rect 41743 2420 42015 2461
rect 42125 2451 42175 2479
rect 42183 2461 42217 2513
rect 42349 2479 42375 2513
rect 42183 2451 42215 2461
rect 42125 2445 42141 2451
rect 42143 2445 42215 2451
rect 42325 2451 42375 2479
rect 42383 2461 42417 2513
rect 42549 2479 42575 2513
rect 42383 2451 42415 2461
rect 42325 2445 42341 2451
rect 42343 2445 42415 2451
rect 42525 2451 42575 2479
rect 42583 2461 42617 2513
rect 42749 2479 42775 2513
rect 42583 2451 42615 2461
rect 42525 2445 42541 2451
rect 42543 2445 42615 2451
rect 42725 2451 42775 2479
rect 42783 2461 42817 2513
rect 42949 2479 42975 2513
rect 42783 2451 42815 2461
rect 42725 2445 42741 2451
rect 42743 2445 42815 2451
rect 42925 2451 42975 2479
rect 42983 2461 43017 2513
rect 43147 2479 43417 2513
rect 43547 2513 45217 2531
rect 43547 2497 43817 2513
rect 42983 2451 43015 2461
rect 42925 2445 42941 2451
rect 42943 2445 43015 2451
rect 43125 2451 43415 2479
rect 43525 2469 43817 2497
rect 43949 2479 43975 2513
rect 43525 2463 43541 2469
rect 43125 2445 43141 2451
rect 41343 2411 41617 2420
rect 39827 2162 39851 2386
rect 39907 2382 39931 2386
rect 39859 2178 39861 2370
rect 39863 2166 39867 2382
rect 39885 2166 39931 2382
rect 39907 2162 39931 2166
rect 39941 2153 40217 2411
rect 40341 2405 40417 2411
rect 40227 2153 40251 2377
rect 40307 2373 40331 2377
rect 40259 2169 40261 2361
rect 40263 2157 40267 2373
rect 40285 2157 40331 2373
rect 40307 2153 40331 2157
rect 40341 2153 40375 2405
rect 39325 2119 39417 2125
rect 39525 2128 39817 2153
rect 39925 2128 40217 2153
rect 39525 2119 39815 2128
rect 39925 2119 39941 2128
rect 39943 2119 40217 2128
rect 40325 2125 40375 2153
rect 40383 2125 40417 2405
rect 40541 2405 40617 2411
rect 40427 2153 40451 2377
rect 40507 2373 40531 2377
rect 40459 2169 40461 2361
rect 40463 2157 40467 2373
rect 40485 2157 40531 2373
rect 40507 2153 40531 2157
rect 40541 2153 40575 2405
rect 40325 2119 40417 2125
rect 40525 2125 40575 2153
rect 40583 2125 40617 2405
rect 40741 2405 40817 2411
rect 40627 2153 40651 2377
rect 40707 2373 40731 2377
rect 40659 2169 40661 2361
rect 40663 2157 40667 2373
rect 40685 2157 40731 2373
rect 40707 2153 40731 2157
rect 40741 2153 40775 2405
rect 40525 2119 40617 2125
rect 40725 2125 40775 2153
rect 40783 2125 40817 2405
rect 40941 2405 41017 2411
rect 40827 2153 40851 2377
rect 40907 2373 40931 2377
rect 40859 2169 40861 2361
rect 40863 2157 40867 2373
rect 40885 2157 40931 2373
rect 40907 2153 40931 2157
rect 40941 2153 40975 2405
rect 40725 2119 40817 2125
rect 40925 2125 40975 2153
rect 40983 2125 41017 2405
rect 41141 2405 41217 2411
rect 41027 2153 41051 2377
rect 41107 2373 41131 2377
rect 41059 2169 41061 2361
rect 41063 2157 41067 2373
rect 41085 2157 41131 2373
rect 41107 2153 41131 2157
rect 41141 2153 41175 2405
rect 40925 2119 41017 2125
rect 41125 2125 41175 2153
rect 41183 2125 41217 2405
rect 41227 2153 41251 2377
rect 41307 2373 41331 2377
rect 41259 2169 41261 2361
rect 41263 2157 41267 2373
rect 41285 2157 41331 2373
rect 41307 2153 41331 2157
rect 41341 2153 41617 2411
rect 41741 2411 42015 2420
rect 42143 2411 42175 2445
rect 42183 2411 42215 2445
rect 42343 2411 42375 2445
rect 42383 2411 42415 2445
rect 42543 2411 42575 2445
rect 42583 2411 42615 2445
rect 42743 2411 42775 2445
rect 42783 2411 42815 2445
rect 42943 2411 42975 2445
rect 42983 2411 43015 2445
rect 43143 2420 43415 2451
rect 43543 2461 43817 2469
rect 43543 2420 43815 2461
rect 43925 2451 43975 2479
rect 43983 2461 44017 2513
rect 44149 2479 44175 2513
rect 43983 2451 44015 2461
rect 43925 2445 43941 2451
rect 43943 2445 44015 2451
rect 44125 2451 44175 2479
rect 44183 2461 44217 2513
rect 44349 2479 44375 2513
rect 44183 2451 44215 2461
rect 44125 2445 44141 2451
rect 44143 2445 44215 2451
rect 44325 2451 44375 2479
rect 44383 2461 44417 2513
rect 44549 2479 44575 2513
rect 44383 2451 44415 2461
rect 44325 2445 44341 2451
rect 44343 2445 44415 2451
rect 44525 2451 44575 2479
rect 44583 2461 44617 2513
rect 44749 2479 44775 2513
rect 44583 2451 44615 2461
rect 44525 2445 44541 2451
rect 44543 2445 44615 2451
rect 44725 2451 44775 2479
rect 44783 2461 44817 2513
rect 44947 2479 45217 2513
rect 45347 2513 47017 2531
rect 45347 2497 45617 2513
rect 44783 2451 44815 2461
rect 44725 2445 44741 2451
rect 44743 2445 44815 2451
rect 44925 2451 45215 2479
rect 45325 2469 45617 2497
rect 45749 2479 45775 2513
rect 45325 2463 45341 2469
rect 44925 2445 44941 2451
rect 43143 2411 43417 2420
rect 41627 2162 41651 2386
rect 41707 2382 41731 2386
rect 41659 2178 41661 2370
rect 41663 2166 41667 2382
rect 41685 2166 41731 2382
rect 41707 2162 41731 2166
rect 41741 2153 42017 2411
rect 42141 2405 42217 2411
rect 42027 2153 42051 2377
rect 42107 2373 42131 2377
rect 42059 2169 42061 2361
rect 42063 2157 42067 2373
rect 42085 2157 42131 2373
rect 42107 2153 42131 2157
rect 42141 2153 42175 2405
rect 41125 2119 41217 2125
rect 41325 2128 41617 2153
rect 41725 2128 42017 2153
rect 41325 2119 41615 2128
rect 41725 2119 41741 2128
rect 41743 2119 42017 2128
rect 42125 2125 42175 2153
rect 42183 2125 42217 2405
rect 42341 2405 42417 2411
rect 42227 2153 42251 2377
rect 42307 2373 42331 2377
rect 42259 2169 42261 2361
rect 42263 2157 42267 2373
rect 42285 2157 42331 2373
rect 42307 2153 42331 2157
rect 42341 2153 42375 2405
rect 42125 2119 42217 2125
rect 42325 2125 42375 2153
rect 42383 2125 42417 2405
rect 42541 2405 42617 2411
rect 42427 2153 42451 2377
rect 42507 2373 42531 2377
rect 42459 2169 42461 2361
rect 42463 2157 42467 2373
rect 42485 2157 42531 2373
rect 42507 2153 42531 2157
rect 42541 2153 42575 2405
rect 42325 2119 42417 2125
rect 42525 2125 42575 2153
rect 42583 2125 42617 2405
rect 42741 2405 42817 2411
rect 42627 2153 42651 2377
rect 42707 2373 42731 2377
rect 42659 2169 42661 2361
rect 42663 2157 42667 2373
rect 42685 2157 42731 2373
rect 42707 2153 42731 2157
rect 42741 2153 42775 2405
rect 42525 2119 42617 2125
rect 42725 2125 42775 2153
rect 42783 2125 42817 2405
rect 42941 2405 43017 2411
rect 42827 2153 42851 2377
rect 42907 2373 42931 2377
rect 42859 2169 42861 2361
rect 42863 2157 42867 2373
rect 42885 2157 42931 2373
rect 42907 2153 42931 2157
rect 42941 2153 42975 2405
rect 42725 2119 42817 2125
rect 42925 2125 42975 2153
rect 42983 2125 43017 2405
rect 43027 2153 43051 2377
rect 43107 2373 43131 2377
rect 43059 2169 43061 2361
rect 43063 2157 43067 2373
rect 43085 2157 43131 2373
rect 43107 2153 43131 2157
rect 43141 2153 43417 2411
rect 43541 2411 43815 2420
rect 43943 2411 43975 2445
rect 43983 2411 44015 2445
rect 44143 2411 44175 2445
rect 44183 2411 44215 2445
rect 44343 2411 44375 2445
rect 44383 2411 44415 2445
rect 44543 2411 44575 2445
rect 44583 2411 44615 2445
rect 44743 2411 44775 2445
rect 44783 2411 44815 2445
rect 44943 2420 45215 2451
rect 45343 2461 45617 2469
rect 45343 2420 45615 2461
rect 45725 2451 45775 2479
rect 45783 2461 45817 2513
rect 45949 2479 45975 2513
rect 45783 2451 45815 2461
rect 45725 2445 45741 2451
rect 45743 2445 45815 2451
rect 45925 2451 45975 2479
rect 45983 2461 46017 2513
rect 46149 2479 46175 2513
rect 45983 2451 46015 2461
rect 45925 2445 45941 2451
rect 45943 2445 46015 2451
rect 46125 2451 46175 2479
rect 46183 2461 46217 2513
rect 46349 2479 46375 2513
rect 46183 2451 46215 2461
rect 46125 2445 46141 2451
rect 46143 2445 46215 2451
rect 46325 2451 46375 2479
rect 46383 2461 46417 2513
rect 46549 2479 46575 2513
rect 46383 2451 46415 2461
rect 46325 2445 46341 2451
rect 46343 2445 46415 2451
rect 46525 2451 46575 2479
rect 46583 2461 46617 2513
rect 46747 2479 47017 2513
rect 47147 2513 48817 2531
rect 47147 2497 47417 2513
rect 46583 2451 46615 2461
rect 46525 2445 46541 2451
rect 46543 2445 46615 2451
rect 46725 2451 47015 2479
rect 47125 2469 47417 2497
rect 47549 2479 47575 2513
rect 47125 2463 47141 2469
rect 46725 2445 46741 2451
rect 44943 2411 45217 2420
rect 43427 2162 43451 2386
rect 43507 2382 43531 2386
rect 43459 2178 43461 2370
rect 43463 2166 43467 2382
rect 43485 2166 43531 2382
rect 43507 2162 43531 2166
rect 43541 2153 43817 2411
rect 43941 2405 44017 2411
rect 43827 2153 43851 2377
rect 43907 2373 43931 2377
rect 43859 2169 43861 2361
rect 43863 2157 43867 2373
rect 43885 2157 43931 2373
rect 43907 2153 43931 2157
rect 43941 2153 43975 2405
rect 42925 2119 43017 2125
rect 43125 2128 43417 2153
rect 43525 2128 43817 2153
rect 43125 2119 43415 2128
rect 43525 2119 43541 2128
rect 43543 2119 43817 2128
rect 43925 2125 43975 2153
rect 43983 2125 44017 2405
rect 44141 2405 44217 2411
rect 44027 2153 44051 2377
rect 44107 2373 44131 2377
rect 44059 2169 44061 2361
rect 44063 2157 44067 2373
rect 44085 2157 44131 2373
rect 44107 2153 44131 2157
rect 44141 2153 44175 2405
rect 43925 2119 44017 2125
rect 44125 2125 44175 2153
rect 44183 2125 44217 2405
rect 44341 2405 44417 2411
rect 44227 2153 44251 2377
rect 44307 2373 44331 2377
rect 44259 2169 44261 2361
rect 44263 2157 44267 2373
rect 44285 2157 44331 2373
rect 44307 2153 44331 2157
rect 44341 2153 44375 2405
rect 44125 2119 44217 2125
rect 44325 2125 44375 2153
rect 44383 2125 44417 2405
rect 44541 2405 44617 2411
rect 44427 2153 44451 2377
rect 44507 2373 44531 2377
rect 44459 2169 44461 2361
rect 44463 2157 44467 2373
rect 44485 2157 44531 2373
rect 44507 2153 44531 2157
rect 44541 2153 44575 2405
rect 44325 2119 44417 2125
rect 44525 2125 44575 2153
rect 44583 2125 44617 2405
rect 44741 2405 44817 2411
rect 44627 2153 44651 2377
rect 44707 2373 44731 2377
rect 44659 2169 44661 2361
rect 44663 2157 44667 2373
rect 44685 2157 44731 2373
rect 44707 2153 44731 2157
rect 44741 2153 44775 2405
rect 44525 2119 44617 2125
rect 44725 2125 44775 2153
rect 44783 2125 44817 2405
rect 44827 2153 44851 2377
rect 44907 2373 44931 2377
rect 44859 2169 44861 2361
rect 44863 2157 44867 2373
rect 44885 2157 44931 2373
rect 44907 2153 44931 2157
rect 44941 2153 45217 2411
rect 45341 2411 45615 2420
rect 45743 2411 45775 2445
rect 45783 2411 45815 2445
rect 45943 2411 45975 2445
rect 45983 2411 46015 2445
rect 46143 2411 46175 2445
rect 46183 2411 46215 2445
rect 46343 2411 46375 2445
rect 46383 2411 46415 2445
rect 46543 2411 46575 2445
rect 46583 2411 46615 2445
rect 46743 2420 47015 2451
rect 47143 2461 47417 2469
rect 47143 2420 47415 2461
rect 47525 2451 47575 2479
rect 47583 2461 47617 2513
rect 47749 2479 47775 2513
rect 47583 2451 47615 2461
rect 47525 2445 47541 2451
rect 47543 2445 47615 2451
rect 47725 2451 47775 2479
rect 47783 2461 47817 2513
rect 47949 2479 47975 2513
rect 47783 2451 47815 2461
rect 47725 2445 47741 2451
rect 47743 2445 47815 2451
rect 47925 2451 47975 2479
rect 47983 2461 48017 2513
rect 48149 2479 48175 2513
rect 47983 2451 48015 2461
rect 47925 2445 47941 2451
rect 47943 2445 48015 2451
rect 48125 2451 48175 2479
rect 48183 2461 48217 2513
rect 48349 2479 48375 2513
rect 48183 2451 48215 2461
rect 48125 2445 48141 2451
rect 48143 2445 48215 2451
rect 48325 2451 48375 2479
rect 48383 2461 48417 2513
rect 48547 2479 48817 2513
rect 48947 2513 50617 2531
rect 48947 2497 49217 2513
rect 48383 2451 48415 2461
rect 48325 2445 48341 2451
rect 48343 2445 48415 2451
rect 48525 2451 48815 2479
rect 48925 2469 49217 2497
rect 49349 2479 49375 2513
rect 48925 2463 48941 2469
rect 48525 2445 48541 2451
rect 46743 2411 47017 2420
rect 45227 2162 45251 2386
rect 45307 2382 45331 2386
rect 45259 2178 45261 2370
rect 45263 2166 45267 2382
rect 45285 2166 45331 2382
rect 45307 2162 45331 2166
rect 45341 2153 45617 2411
rect 45741 2405 45817 2411
rect 45627 2153 45651 2377
rect 45707 2373 45731 2377
rect 45659 2169 45661 2361
rect 45663 2157 45667 2373
rect 45685 2157 45731 2373
rect 45707 2153 45731 2157
rect 45741 2153 45775 2405
rect 44725 2119 44817 2125
rect 44925 2128 45217 2153
rect 45325 2128 45617 2153
rect 44925 2119 45215 2128
rect 45325 2119 45341 2128
rect 45343 2119 45617 2128
rect 45725 2125 45775 2153
rect 45783 2125 45817 2405
rect 45941 2405 46017 2411
rect 45827 2153 45851 2377
rect 45907 2373 45931 2377
rect 45859 2169 45861 2361
rect 45863 2157 45867 2373
rect 45885 2157 45931 2373
rect 45907 2153 45931 2157
rect 45941 2153 45975 2405
rect 45725 2119 45817 2125
rect 45925 2125 45975 2153
rect 45983 2125 46017 2405
rect 46141 2405 46217 2411
rect 46027 2153 46051 2377
rect 46107 2373 46131 2377
rect 46059 2169 46061 2361
rect 46063 2157 46067 2373
rect 46085 2157 46131 2373
rect 46107 2153 46131 2157
rect 46141 2153 46175 2405
rect 45925 2119 46017 2125
rect 46125 2125 46175 2153
rect 46183 2125 46217 2405
rect 46341 2405 46417 2411
rect 46227 2153 46251 2377
rect 46307 2373 46331 2377
rect 46259 2169 46261 2361
rect 46263 2157 46267 2373
rect 46285 2157 46331 2373
rect 46307 2153 46331 2157
rect 46341 2153 46375 2405
rect 46125 2119 46217 2125
rect 46325 2125 46375 2153
rect 46383 2125 46417 2405
rect 46541 2405 46617 2411
rect 46427 2153 46451 2377
rect 46507 2373 46531 2377
rect 46459 2169 46461 2361
rect 46463 2157 46467 2373
rect 46485 2157 46531 2373
rect 46507 2153 46531 2157
rect 46541 2153 46575 2405
rect 46325 2119 46417 2125
rect 46525 2125 46575 2153
rect 46583 2125 46617 2405
rect 46627 2153 46651 2377
rect 46707 2373 46731 2377
rect 46659 2169 46661 2361
rect 46663 2157 46667 2373
rect 46685 2157 46731 2373
rect 46707 2153 46731 2157
rect 46741 2153 47017 2411
rect 47141 2411 47415 2420
rect 47543 2411 47575 2445
rect 47583 2411 47615 2445
rect 47743 2411 47775 2445
rect 47783 2411 47815 2445
rect 47943 2411 47975 2445
rect 47983 2411 48015 2445
rect 48143 2411 48175 2445
rect 48183 2411 48215 2445
rect 48343 2411 48375 2445
rect 48383 2411 48415 2445
rect 48543 2420 48815 2451
rect 48943 2461 49217 2469
rect 48943 2420 49215 2461
rect 49325 2451 49375 2479
rect 49383 2461 49417 2513
rect 49549 2479 49575 2513
rect 49383 2451 49415 2461
rect 49325 2445 49341 2451
rect 49343 2445 49415 2451
rect 49525 2451 49575 2479
rect 49583 2461 49617 2513
rect 49749 2479 49775 2513
rect 49583 2451 49615 2461
rect 49525 2445 49541 2451
rect 49543 2445 49615 2451
rect 49725 2451 49775 2479
rect 49783 2461 49817 2513
rect 49949 2479 49975 2513
rect 49783 2451 49815 2461
rect 49725 2445 49741 2451
rect 49743 2445 49815 2451
rect 49925 2451 49975 2479
rect 49983 2461 50017 2513
rect 50149 2479 50175 2513
rect 49983 2451 50015 2461
rect 49925 2445 49941 2451
rect 49943 2445 50015 2451
rect 50125 2451 50175 2479
rect 50183 2461 50217 2513
rect 50347 2479 50617 2513
rect 50747 2513 52417 2531
rect 50747 2497 51017 2513
rect 50183 2451 50215 2461
rect 50125 2445 50141 2451
rect 50143 2445 50215 2451
rect 50325 2451 50615 2479
rect 50725 2469 51017 2497
rect 51149 2479 51175 2513
rect 50725 2463 50741 2469
rect 50325 2445 50341 2451
rect 48543 2411 48817 2420
rect 47027 2162 47051 2386
rect 47107 2382 47131 2386
rect 47059 2178 47061 2370
rect 47063 2166 47067 2382
rect 47085 2166 47131 2382
rect 47107 2162 47131 2166
rect 47141 2153 47417 2411
rect 47541 2405 47617 2411
rect 47427 2153 47451 2377
rect 47507 2373 47531 2377
rect 47459 2169 47461 2361
rect 47463 2157 47467 2373
rect 47485 2157 47531 2373
rect 47507 2153 47531 2157
rect 47541 2153 47575 2405
rect 46525 2119 46617 2125
rect 46725 2128 47017 2153
rect 47125 2128 47417 2153
rect 46725 2119 47015 2128
rect 47125 2119 47141 2128
rect 47143 2119 47417 2128
rect 47525 2125 47575 2153
rect 47583 2125 47617 2405
rect 47741 2405 47817 2411
rect 47627 2153 47651 2377
rect 47707 2373 47731 2377
rect 47659 2169 47661 2361
rect 47663 2157 47667 2373
rect 47685 2157 47731 2373
rect 47707 2153 47731 2157
rect 47741 2153 47775 2405
rect 47525 2119 47617 2125
rect 47725 2125 47775 2153
rect 47783 2125 47817 2405
rect 47941 2405 48017 2411
rect 47827 2153 47851 2377
rect 47907 2373 47931 2377
rect 47859 2169 47861 2361
rect 47863 2157 47867 2373
rect 47885 2157 47931 2373
rect 47907 2153 47931 2157
rect 47941 2153 47975 2405
rect 47725 2119 47817 2125
rect 47925 2125 47975 2153
rect 47983 2125 48017 2405
rect 48141 2405 48217 2411
rect 48027 2153 48051 2377
rect 48107 2373 48131 2377
rect 48059 2169 48061 2361
rect 48063 2157 48067 2373
rect 48085 2157 48131 2373
rect 48107 2153 48131 2157
rect 48141 2153 48175 2405
rect 47925 2119 48017 2125
rect 48125 2125 48175 2153
rect 48183 2125 48217 2405
rect 48341 2405 48417 2411
rect 48227 2153 48251 2377
rect 48307 2373 48331 2377
rect 48259 2169 48261 2361
rect 48263 2157 48267 2373
rect 48285 2157 48331 2373
rect 48307 2153 48331 2157
rect 48341 2153 48375 2405
rect 48125 2119 48217 2125
rect 48325 2125 48375 2153
rect 48383 2125 48417 2405
rect 48427 2153 48451 2377
rect 48507 2373 48531 2377
rect 48459 2169 48461 2361
rect 48463 2157 48467 2373
rect 48485 2157 48531 2373
rect 48507 2153 48531 2157
rect 48541 2153 48817 2411
rect 48941 2411 49215 2420
rect 49343 2411 49375 2445
rect 49383 2411 49415 2445
rect 49543 2411 49575 2445
rect 49583 2411 49615 2445
rect 49743 2411 49775 2445
rect 49783 2411 49815 2445
rect 49943 2411 49975 2445
rect 49983 2411 50015 2445
rect 50143 2411 50175 2445
rect 50183 2411 50215 2445
rect 50343 2420 50615 2451
rect 50743 2461 51017 2469
rect 50743 2420 51015 2461
rect 51125 2451 51175 2479
rect 51183 2461 51217 2513
rect 51349 2479 51375 2513
rect 51183 2451 51215 2461
rect 51125 2445 51141 2451
rect 51143 2445 51215 2451
rect 51325 2451 51375 2479
rect 51383 2461 51417 2513
rect 51549 2479 51575 2513
rect 51383 2451 51415 2461
rect 51325 2445 51341 2451
rect 51343 2445 51415 2451
rect 51525 2451 51575 2479
rect 51583 2461 51617 2513
rect 51749 2479 51775 2513
rect 51583 2451 51615 2461
rect 51525 2445 51541 2451
rect 51543 2445 51615 2451
rect 51725 2451 51775 2479
rect 51783 2461 51817 2513
rect 51949 2479 51975 2513
rect 51783 2451 51815 2461
rect 51725 2445 51741 2451
rect 51743 2445 51815 2451
rect 51925 2451 51975 2479
rect 51983 2461 52017 2513
rect 52147 2479 52417 2513
rect 52547 2513 54217 2531
rect 52547 2497 52817 2513
rect 51983 2451 52015 2461
rect 51925 2445 51941 2451
rect 51943 2445 52015 2451
rect 52125 2451 52415 2479
rect 52525 2469 52817 2497
rect 52949 2479 52975 2513
rect 52525 2463 52541 2469
rect 52125 2445 52141 2451
rect 50343 2411 50617 2420
rect 48827 2162 48851 2386
rect 48907 2382 48931 2386
rect 48859 2178 48861 2370
rect 48863 2166 48867 2382
rect 48885 2166 48931 2382
rect 48907 2162 48931 2166
rect 48941 2153 49217 2411
rect 49341 2405 49417 2411
rect 49227 2153 49251 2377
rect 49307 2373 49331 2377
rect 49259 2169 49261 2361
rect 49263 2157 49267 2373
rect 49285 2157 49331 2373
rect 49307 2153 49331 2157
rect 49341 2153 49375 2405
rect 48325 2119 48417 2125
rect 48525 2128 48817 2153
rect 48925 2128 49217 2153
rect 48525 2119 48815 2128
rect 48925 2119 48941 2128
rect 48943 2119 49217 2128
rect 49325 2125 49375 2153
rect 49383 2125 49417 2405
rect 49541 2405 49617 2411
rect 49427 2153 49451 2377
rect 49507 2373 49531 2377
rect 49459 2169 49461 2361
rect 49463 2157 49467 2373
rect 49485 2157 49531 2373
rect 49507 2153 49531 2157
rect 49541 2153 49575 2405
rect 49325 2119 49417 2125
rect 49525 2125 49575 2153
rect 49583 2125 49617 2405
rect 49741 2405 49817 2411
rect 49627 2153 49651 2377
rect 49707 2373 49731 2377
rect 49659 2169 49661 2361
rect 49663 2157 49667 2373
rect 49685 2157 49731 2373
rect 49707 2153 49731 2157
rect 49741 2153 49775 2405
rect 49525 2119 49617 2125
rect 49725 2125 49775 2153
rect 49783 2125 49817 2405
rect 49941 2405 50017 2411
rect 49827 2153 49851 2377
rect 49907 2373 49931 2377
rect 49859 2169 49861 2361
rect 49863 2157 49867 2373
rect 49885 2157 49931 2373
rect 49907 2153 49931 2157
rect 49941 2153 49975 2405
rect 49725 2119 49817 2125
rect 49925 2125 49975 2153
rect 49983 2125 50017 2405
rect 50141 2405 50217 2411
rect 50027 2153 50051 2377
rect 50107 2373 50131 2377
rect 50059 2169 50061 2361
rect 50063 2157 50067 2373
rect 50085 2157 50131 2373
rect 50107 2153 50131 2157
rect 50141 2153 50175 2405
rect 49925 2119 50017 2125
rect 50125 2125 50175 2153
rect 50183 2125 50217 2405
rect 50227 2153 50251 2377
rect 50307 2373 50331 2377
rect 50259 2169 50261 2361
rect 50263 2157 50267 2373
rect 50285 2157 50331 2373
rect 50307 2153 50331 2157
rect 50341 2153 50617 2411
rect 50741 2411 51015 2420
rect 51143 2411 51175 2445
rect 51183 2411 51215 2445
rect 51343 2411 51375 2445
rect 51383 2411 51415 2445
rect 51543 2411 51575 2445
rect 51583 2411 51615 2445
rect 51743 2411 51775 2445
rect 51783 2411 51815 2445
rect 51943 2411 51975 2445
rect 51983 2411 52015 2445
rect 52143 2420 52415 2451
rect 52543 2461 52817 2469
rect 52543 2420 52815 2461
rect 52925 2451 52975 2479
rect 52983 2461 53017 2513
rect 53149 2479 53175 2513
rect 52983 2451 53015 2461
rect 52925 2445 52941 2451
rect 52943 2445 53015 2451
rect 53125 2451 53175 2479
rect 53183 2461 53217 2513
rect 53349 2479 53375 2513
rect 53183 2451 53215 2461
rect 53125 2445 53141 2451
rect 53143 2445 53215 2451
rect 53325 2451 53375 2479
rect 53383 2461 53417 2513
rect 53549 2479 53575 2513
rect 53383 2451 53415 2461
rect 53325 2445 53341 2451
rect 53343 2445 53415 2451
rect 53525 2451 53575 2479
rect 53583 2461 53617 2513
rect 53749 2479 53775 2513
rect 53583 2451 53615 2461
rect 53525 2445 53541 2451
rect 53543 2445 53615 2451
rect 53725 2451 53775 2479
rect 53783 2461 53817 2513
rect 53947 2479 54217 2513
rect 54347 2513 56017 2531
rect 54347 2497 54617 2513
rect 53783 2451 53815 2461
rect 53725 2445 53741 2451
rect 53743 2445 53815 2451
rect 53925 2451 54215 2479
rect 54325 2469 54617 2497
rect 54749 2479 54775 2513
rect 54325 2463 54341 2469
rect 53925 2445 53941 2451
rect 52143 2411 52417 2420
rect 50627 2162 50651 2386
rect 50707 2382 50731 2386
rect 50659 2178 50661 2370
rect 50663 2166 50667 2382
rect 50685 2166 50731 2382
rect 50707 2162 50731 2166
rect 50741 2153 51017 2411
rect 51141 2405 51217 2411
rect 51027 2153 51051 2377
rect 51107 2373 51131 2377
rect 51059 2169 51061 2361
rect 51063 2157 51067 2373
rect 51085 2157 51131 2373
rect 51107 2153 51131 2157
rect 51141 2153 51175 2405
rect 50125 2119 50217 2125
rect 50325 2128 50617 2153
rect 50725 2128 51017 2153
rect 50325 2119 50615 2128
rect 50725 2119 50741 2128
rect 50743 2119 51017 2128
rect 51125 2125 51175 2153
rect 51183 2125 51217 2405
rect 51341 2405 51417 2411
rect 51227 2153 51251 2377
rect 51307 2373 51331 2377
rect 51259 2169 51261 2361
rect 51263 2157 51267 2373
rect 51285 2157 51331 2373
rect 51307 2153 51331 2157
rect 51341 2153 51375 2405
rect 51125 2119 51217 2125
rect 51325 2125 51375 2153
rect 51383 2125 51417 2405
rect 51541 2405 51617 2411
rect 51427 2153 51451 2377
rect 51507 2373 51531 2377
rect 51459 2169 51461 2361
rect 51463 2157 51467 2373
rect 51485 2157 51531 2373
rect 51507 2153 51531 2157
rect 51541 2153 51575 2405
rect 51325 2119 51417 2125
rect 51525 2125 51575 2153
rect 51583 2125 51617 2405
rect 51741 2405 51817 2411
rect 51627 2153 51651 2377
rect 51707 2373 51731 2377
rect 51659 2169 51661 2361
rect 51663 2157 51667 2373
rect 51685 2157 51731 2373
rect 51707 2153 51731 2157
rect 51741 2153 51775 2405
rect 51525 2119 51617 2125
rect 51725 2125 51775 2153
rect 51783 2125 51817 2405
rect 51941 2405 52017 2411
rect 51827 2153 51851 2377
rect 51907 2373 51931 2377
rect 51859 2169 51861 2361
rect 51863 2157 51867 2373
rect 51885 2157 51931 2373
rect 51907 2153 51931 2157
rect 51941 2153 51975 2405
rect 51725 2119 51817 2125
rect 51925 2125 51975 2153
rect 51983 2125 52017 2405
rect 52027 2153 52051 2377
rect 52107 2373 52131 2377
rect 52059 2169 52061 2361
rect 52063 2157 52067 2373
rect 52085 2157 52131 2373
rect 52107 2153 52131 2157
rect 52141 2153 52417 2411
rect 52541 2411 52815 2420
rect 52943 2411 52975 2445
rect 52983 2411 53015 2445
rect 53143 2411 53175 2445
rect 53183 2411 53215 2445
rect 53343 2411 53375 2445
rect 53383 2411 53415 2445
rect 53543 2411 53575 2445
rect 53583 2411 53615 2445
rect 53743 2411 53775 2445
rect 53783 2411 53815 2445
rect 53943 2420 54215 2451
rect 54343 2461 54617 2469
rect 54343 2420 54615 2461
rect 54725 2451 54775 2479
rect 54783 2461 54817 2513
rect 54949 2479 54975 2513
rect 54783 2451 54815 2461
rect 54725 2445 54741 2451
rect 54743 2445 54815 2451
rect 54925 2451 54975 2479
rect 54983 2461 55017 2513
rect 55149 2479 55175 2513
rect 54983 2451 55015 2461
rect 54925 2445 54941 2451
rect 54943 2445 55015 2451
rect 55125 2451 55175 2479
rect 55183 2461 55217 2513
rect 55349 2479 55375 2513
rect 55183 2451 55215 2461
rect 55125 2445 55141 2451
rect 55143 2445 55215 2451
rect 55325 2451 55375 2479
rect 55383 2461 55417 2513
rect 55549 2479 55575 2513
rect 55383 2451 55415 2461
rect 55325 2445 55341 2451
rect 55343 2445 55415 2451
rect 55525 2451 55575 2479
rect 55583 2461 55617 2513
rect 55747 2479 56017 2513
rect 56147 2513 57817 2531
rect 56147 2497 56417 2513
rect 55583 2451 55615 2461
rect 55525 2445 55541 2451
rect 55543 2445 55615 2451
rect 55725 2451 56015 2479
rect 56125 2469 56417 2497
rect 56549 2479 56575 2513
rect 56125 2463 56141 2469
rect 55725 2445 55741 2451
rect 53943 2411 54217 2420
rect 52427 2162 52451 2386
rect 52507 2382 52531 2386
rect 52459 2178 52461 2370
rect 52463 2166 52467 2382
rect 52485 2166 52531 2382
rect 52507 2162 52531 2166
rect 52541 2153 52817 2411
rect 52941 2405 53017 2411
rect 52827 2153 52851 2377
rect 52907 2373 52931 2377
rect 52859 2169 52861 2361
rect 52863 2157 52867 2373
rect 52885 2157 52931 2373
rect 52907 2153 52931 2157
rect 52941 2153 52975 2405
rect 51925 2119 52017 2125
rect 52125 2128 52417 2153
rect 52525 2128 52817 2153
rect 52125 2119 52415 2128
rect 52525 2119 52541 2128
rect 52543 2119 52817 2128
rect 52925 2125 52975 2153
rect 52983 2125 53017 2405
rect 53141 2405 53217 2411
rect 53027 2153 53051 2377
rect 53107 2373 53131 2377
rect 53059 2169 53061 2361
rect 53063 2157 53067 2373
rect 53085 2157 53131 2373
rect 53107 2153 53131 2157
rect 53141 2153 53175 2405
rect 52925 2119 53017 2125
rect 53125 2125 53175 2153
rect 53183 2125 53217 2405
rect 53341 2405 53417 2411
rect 53227 2153 53251 2377
rect 53307 2373 53331 2377
rect 53259 2169 53261 2361
rect 53263 2157 53267 2373
rect 53285 2157 53331 2373
rect 53307 2153 53331 2157
rect 53341 2153 53375 2405
rect 53125 2119 53217 2125
rect 53325 2125 53375 2153
rect 53383 2125 53417 2405
rect 53541 2405 53617 2411
rect 53427 2153 53451 2377
rect 53507 2373 53531 2377
rect 53459 2169 53461 2361
rect 53463 2157 53467 2373
rect 53485 2157 53531 2373
rect 53507 2153 53531 2157
rect 53541 2153 53575 2405
rect 53325 2119 53417 2125
rect 53525 2125 53575 2153
rect 53583 2125 53617 2405
rect 53741 2405 53817 2411
rect 53627 2153 53651 2377
rect 53707 2373 53731 2377
rect 53659 2169 53661 2361
rect 53663 2157 53667 2373
rect 53685 2157 53731 2373
rect 53707 2153 53731 2157
rect 53741 2153 53775 2405
rect 53525 2119 53617 2125
rect 53725 2125 53775 2153
rect 53783 2125 53817 2405
rect 53827 2153 53851 2377
rect 53907 2373 53931 2377
rect 53859 2169 53861 2361
rect 53863 2157 53867 2373
rect 53885 2157 53931 2373
rect 53907 2153 53931 2157
rect 53941 2153 54217 2411
rect 54341 2411 54615 2420
rect 54743 2411 54775 2445
rect 54783 2411 54815 2445
rect 54943 2411 54975 2445
rect 54983 2411 55015 2445
rect 55143 2411 55175 2445
rect 55183 2411 55215 2445
rect 55343 2411 55375 2445
rect 55383 2411 55415 2445
rect 55543 2411 55575 2445
rect 55583 2411 55615 2445
rect 55743 2420 56015 2451
rect 56143 2461 56417 2469
rect 56143 2420 56415 2461
rect 56525 2451 56575 2479
rect 56583 2461 56617 2513
rect 56749 2479 56775 2513
rect 56583 2451 56615 2461
rect 56525 2445 56541 2451
rect 56543 2445 56615 2451
rect 56725 2451 56775 2479
rect 56783 2461 56817 2513
rect 56949 2479 56975 2513
rect 56783 2451 56815 2461
rect 56725 2445 56741 2451
rect 56743 2445 56815 2451
rect 56925 2451 56975 2479
rect 56983 2461 57017 2513
rect 57149 2479 57175 2513
rect 56983 2451 57015 2461
rect 56925 2445 56941 2451
rect 56943 2445 57015 2451
rect 57125 2451 57175 2479
rect 57183 2461 57217 2513
rect 57349 2479 57375 2513
rect 57183 2451 57215 2461
rect 57125 2445 57141 2451
rect 57143 2445 57215 2451
rect 57325 2451 57375 2479
rect 57383 2461 57417 2513
rect 57547 2479 57817 2513
rect 57947 2513 59617 2531
rect 57947 2497 58217 2513
rect 57383 2451 57415 2461
rect 57325 2445 57341 2451
rect 57343 2445 57415 2451
rect 57525 2451 57815 2479
rect 57925 2469 58217 2497
rect 58349 2479 58375 2513
rect 57925 2463 57941 2469
rect 57525 2445 57541 2451
rect 55743 2411 56017 2420
rect 54227 2162 54251 2386
rect 54307 2382 54331 2386
rect 54259 2178 54261 2370
rect 54263 2166 54267 2382
rect 54285 2166 54331 2382
rect 54307 2162 54331 2166
rect 54341 2153 54617 2411
rect 54741 2405 54817 2411
rect 54627 2153 54651 2377
rect 54707 2373 54731 2377
rect 54659 2169 54661 2361
rect 54663 2157 54667 2373
rect 54685 2157 54731 2373
rect 54707 2153 54731 2157
rect 54741 2153 54775 2405
rect 53725 2119 53817 2125
rect 53925 2128 54217 2153
rect 54325 2128 54617 2153
rect 53925 2119 54215 2128
rect 54325 2119 54341 2128
rect 54343 2119 54617 2128
rect 54725 2125 54775 2153
rect 54783 2125 54817 2405
rect 54941 2405 55017 2411
rect 54827 2153 54851 2377
rect 54907 2373 54931 2377
rect 54859 2169 54861 2361
rect 54863 2157 54867 2373
rect 54885 2157 54931 2373
rect 54907 2153 54931 2157
rect 54941 2153 54975 2405
rect 54725 2119 54817 2125
rect 54925 2125 54975 2153
rect 54983 2125 55017 2405
rect 55141 2405 55217 2411
rect 55027 2153 55051 2377
rect 55107 2373 55131 2377
rect 55059 2169 55061 2361
rect 55063 2157 55067 2373
rect 55085 2157 55131 2373
rect 55107 2153 55131 2157
rect 55141 2153 55175 2405
rect 54925 2119 55017 2125
rect 55125 2125 55175 2153
rect 55183 2125 55217 2405
rect 55341 2405 55417 2411
rect 55227 2153 55251 2377
rect 55307 2373 55331 2377
rect 55259 2169 55261 2361
rect 55263 2157 55267 2373
rect 55285 2157 55331 2373
rect 55307 2153 55331 2157
rect 55341 2153 55375 2405
rect 55125 2119 55217 2125
rect 55325 2125 55375 2153
rect 55383 2125 55417 2405
rect 55541 2405 55617 2411
rect 55427 2153 55451 2377
rect 55507 2373 55531 2377
rect 55459 2169 55461 2361
rect 55463 2157 55467 2373
rect 55485 2157 55531 2373
rect 55507 2153 55531 2157
rect 55541 2153 55575 2405
rect 55325 2119 55417 2125
rect 55525 2125 55575 2153
rect 55583 2125 55617 2405
rect 55627 2153 55651 2377
rect 55707 2373 55731 2377
rect 55659 2169 55661 2361
rect 55663 2157 55667 2373
rect 55685 2157 55731 2373
rect 55707 2153 55731 2157
rect 55741 2153 56017 2411
rect 56141 2411 56415 2420
rect 56543 2411 56575 2445
rect 56583 2411 56615 2445
rect 56743 2411 56775 2445
rect 56783 2411 56815 2445
rect 56943 2411 56975 2445
rect 56983 2411 57015 2445
rect 57143 2411 57175 2445
rect 57183 2411 57215 2445
rect 57343 2411 57375 2445
rect 57383 2411 57415 2445
rect 57543 2420 57815 2451
rect 57943 2461 58217 2469
rect 57943 2420 58215 2461
rect 58325 2451 58375 2479
rect 58383 2461 58417 2513
rect 58549 2479 58575 2513
rect 58383 2451 58415 2461
rect 58325 2445 58341 2451
rect 58343 2445 58415 2451
rect 58525 2451 58575 2479
rect 58583 2461 58617 2513
rect 58749 2479 58775 2513
rect 58583 2451 58615 2461
rect 58525 2445 58541 2451
rect 58543 2445 58615 2451
rect 58725 2451 58775 2479
rect 58783 2461 58817 2513
rect 58949 2479 58975 2513
rect 58783 2451 58815 2461
rect 58725 2445 58741 2451
rect 58743 2445 58815 2451
rect 58925 2451 58975 2479
rect 58983 2461 59017 2513
rect 59149 2479 59175 2513
rect 58983 2451 59015 2461
rect 58925 2445 58941 2451
rect 58943 2445 59015 2451
rect 59125 2451 59175 2479
rect 59183 2461 59217 2513
rect 59347 2479 59617 2513
rect 59747 2513 61417 2531
rect 59747 2497 60017 2513
rect 59183 2451 59215 2461
rect 59125 2445 59141 2451
rect 59143 2445 59215 2451
rect 59325 2451 59615 2479
rect 59725 2469 60017 2497
rect 60149 2479 60175 2513
rect 59725 2463 59741 2469
rect 59325 2445 59341 2451
rect 57543 2411 57817 2420
rect 56027 2162 56051 2386
rect 56107 2382 56131 2386
rect 56059 2178 56061 2370
rect 56063 2166 56067 2382
rect 56085 2166 56131 2382
rect 56107 2162 56131 2166
rect 56141 2153 56417 2411
rect 56541 2405 56617 2411
rect 56427 2153 56451 2377
rect 56507 2373 56531 2377
rect 56459 2169 56461 2361
rect 56463 2157 56467 2373
rect 56485 2157 56531 2373
rect 56507 2153 56531 2157
rect 56541 2153 56575 2405
rect 55525 2119 55617 2125
rect 55725 2128 56017 2153
rect 56125 2128 56417 2153
rect 55725 2119 56015 2128
rect 56125 2119 56141 2128
rect 56143 2119 56417 2128
rect 56525 2125 56575 2153
rect 56583 2125 56617 2405
rect 56741 2405 56817 2411
rect 56627 2153 56651 2377
rect 56707 2373 56731 2377
rect 56659 2169 56661 2361
rect 56663 2157 56667 2373
rect 56685 2157 56731 2373
rect 56707 2153 56731 2157
rect 56741 2153 56775 2405
rect 56525 2119 56617 2125
rect 56725 2125 56775 2153
rect 56783 2125 56817 2405
rect 56941 2405 57017 2411
rect 56827 2153 56851 2377
rect 56907 2373 56931 2377
rect 56859 2169 56861 2361
rect 56863 2157 56867 2373
rect 56885 2157 56931 2373
rect 56907 2153 56931 2157
rect 56941 2153 56975 2405
rect 56725 2119 56817 2125
rect 56925 2125 56975 2153
rect 56983 2125 57017 2405
rect 57141 2405 57217 2411
rect 57027 2153 57051 2377
rect 57107 2373 57131 2377
rect 57059 2169 57061 2361
rect 57063 2157 57067 2373
rect 57085 2157 57131 2373
rect 57107 2153 57131 2157
rect 57141 2153 57175 2405
rect 56925 2119 57017 2125
rect 57125 2125 57175 2153
rect 57183 2125 57217 2405
rect 57341 2405 57417 2411
rect 57227 2153 57251 2377
rect 57307 2373 57331 2377
rect 57259 2169 57261 2361
rect 57263 2157 57267 2373
rect 57285 2157 57331 2373
rect 57307 2153 57331 2157
rect 57341 2153 57375 2405
rect 57125 2119 57217 2125
rect 57325 2125 57375 2153
rect 57383 2125 57417 2405
rect 57427 2153 57451 2377
rect 57507 2373 57531 2377
rect 57459 2169 57461 2361
rect 57463 2157 57467 2373
rect 57485 2157 57531 2373
rect 57507 2153 57531 2157
rect 57541 2153 57817 2411
rect 57941 2411 58215 2420
rect 58343 2411 58375 2445
rect 58383 2411 58415 2445
rect 58543 2411 58575 2445
rect 58583 2411 58615 2445
rect 58743 2411 58775 2445
rect 58783 2411 58815 2445
rect 58943 2411 58975 2445
rect 58983 2411 59015 2445
rect 59143 2411 59175 2445
rect 59183 2411 59215 2445
rect 59343 2420 59615 2451
rect 59743 2461 60017 2469
rect 59743 2420 60015 2461
rect 60125 2451 60175 2479
rect 60183 2461 60217 2513
rect 60349 2479 60375 2513
rect 60183 2451 60215 2461
rect 60125 2445 60141 2451
rect 60143 2445 60215 2451
rect 60325 2451 60375 2479
rect 60383 2461 60417 2513
rect 60549 2479 60575 2513
rect 60383 2451 60415 2461
rect 60325 2445 60341 2451
rect 60343 2445 60415 2451
rect 60525 2451 60575 2479
rect 60583 2461 60617 2513
rect 60749 2479 60775 2513
rect 60583 2451 60615 2461
rect 60525 2445 60541 2451
rect 60543 2445 60615 2451
rect 60725 2451 60775 2479
rect 60783 2461 60817 2513
rect 60949 2479 60975 2513
rect 60783 2451 60815 2461
rect 60725 2445 60741 2451
rect 60743 2445 60815 2451
rect 60925 2451 60975 2479
rect 60983 2461 61017 2513
rect 61147 2479 61417 2513
rect 61547 2513 63217 2531
rect 61547 2497 61817 2513
rect 60983 2451 61015 2461
rect 60925 2445 60941 2451
rect 60943 2445 61015 2451
rect 61125 2451 61415 2479
rect 61525 2469 61817 2497
rect 61949 2479 61975 2513
rect 61525 2463 61541 2469
rect 61125 2445 61141 2451
rect 59343 2411 59617 2420
rect 57827 2162 57851 2386
rect 57907 2382 57931 2386
rect 57859 2178 57861 2370
rect 57863 2166 57867 2382
rect 57885 2166 57931 2382
rect 57907 2162 57931 2166
rect 57941 2153 58217 2411
rect 58341 2405 58417 2411
rect 58227 2153 58251 2377
rect 58307 2373 58331 2377
rect 58259 2169 58261 2361
rect 58263 2157 58267 2373
rect 58285 2157 58331 2373
rect 58307 2153 58331 2157
rect 58341 2153 58375 2405
rect 57325 2119 57417 2125
rect 57525 2128 57817 2153
rect 57925 2128 58217 2153
rect 57525 2119 57815 2128
rect 57925 2119 57941 2128
rect 57943 2119 58217 2128
rect 58325 2125 58375 2153
rect 58383 2125 58417 2405
rect 58541 2405 58617 2411
rect 58427 2153 58451 2377
rect 58507 2373 58531 2377
rect 58459 2169 58461 2361
rect 58463 2157 58467 2373
rect 58485 2157 58531 2373
rect 58507 2153 58531 2157
rect 58541 2153 58575 2405
rect 58325 2119 58417 2125
rect 58525 2125 58575 2153
rect 58583 2125 58617 2405
rect 58741 2405 58817 2411
rect 58627 2153 58651 2377
rect 58707 2373 58731 2377
rect 58659 2169 58661 2361
rect 58663 2157 58667 2373
rect 58685 2157 58731 2373
rect 58707 2153 58731 2157
rect 58741 2153 58775 2405
rect 58525 2119 58617 2125
rect 58725 2125 58775 2153
rect 58783 2125 58817 2405
rect 58941 2405 59017 2411
rect 58827 2153 58851 2377
rect 58907 2373 58931 2377
rect 58859 2169 58861 2361
rect 58863 2157 58867 2373
rect 58885 2157 58931 2373
rect 58907 2153 58931 2157
rect 58941 2153 58975 2405
rect 58725 2119 58817 2125
rect 58925 2125 58975 2153
rect 58983 2125 59017 2405
rect 59141 2405 59217 2411
rect 59027 2153 59051 2377
rect 59107 2373 59131 2377
rect 59059 2169 59061 2361
rect 59063 2157 59067 2373
rect 59085 2157 59131 2373
rect 59107 2153 59131 2157
rect 59141 2153 59175 2405
rect 58925 2119 59017 2125
rect 59125 2125 59175 2153
rect 59183 2125 59217 2405
rect 59227 2153 59251 2377
rect 59307 2373 59331 2377
rect 59259 2169 59261 2361
rect 59263 2157 59267 2373
rect 59285 2157 59331 2373
rect 59307 2153 59331 2157
rect 59341 2153 59617 2411
rect 59741 2411 60015 2420
rect 60143 2411 60175 2445
rect 60183 2411 60215 2445
rect 60343 2411 60375 2445
rect 60383 2411 60415 2445
rect 60543 2411 60575 2445
rect 60583 2411 60615 2445
rect 60743 2411 60775 2445
rect 60783 2411 60815 2445
rect 60943 2411 60975 2445
rect 60983 2411 61015 2445
rect 61143 2420 61415 2451
rect 61543 2461 61817 2469
rect 61543 2420 61815 2461
rect 61925 2451 61975 2479
rect 61983 2461 62017 2513
rect 62149 2479 62175 2513
rect 61983 2451 62015 2461
rect 61925 2445 61941 2451
rect 61943 2445 62015 2451
rect 62125 2451 62175 2479
rect 62183 2461 62217 2513
rect 62349 2479 62375 2513
rect 62183 2451 62215 2461
rect 62125 2445 62141 2451
rect 62143 2445 62215 2451
rect 62325 2451 62375 2479
rect 62383 2461 62417 2513
rect 62549 2479 62575 2513
rect 62383 2451 62415 2461
rect 62325 2445 62341 2451
rect 62343 2445 62415 2451
rect 62525 2451 62575 2479
rect 62583 2461 62617 2513
rect 62749 2479 62775 2513
rect 62583 2451 62615 2461
rect 62525 2445 62541 2451
rect 62543 2445 62615 2451
rect 62725 2451 62775 2479
rect 62783 2461 62817 2513
rect 62947 2479 63217 2513
rect 63347 2513 65017 2531
rect 63347 2497 63617 2513
rect 62783 2451 62815 2461
rect 62725 2445 62741 2451
rect 62743 2445 62815 2451
rect 62925 2451 63215 2479
rect 63325 2469 63617 2497
rect 63749 2479 63775 2513
rect 63325 2463 63341 2469
rect 62925 2445 62941 2451
rect 61143 2411 61417 2420
rect 59627 2162 59651 2386
rect 59707 2382 59731 2386
rect 59659 2178 59661 2370
rect 59663 2166 59667 2382
rect 59685 2166 59731 2382
rect 59707 2162 59731 2166
rect 59741 2153 60017 2411
rect 60141 2405 60217 2411
rect 60027 2153 60051 2377
rect 60107 2373 60131 2377
rect 60059 2169 60061 2361
rect 60063 2157 60067 2373
rect 60085 2157 60131 2373
rect 60107 2153 60131 2157
rect 60141 2153 60175 2405
rect 59125 2119 59217 2125
rect 59325 2128 59617 2153
rect 59725 2128 60017 2153
rect 59325 2119 59615 2128
rect 59725 2119 59741 2128
rect 59743 2119 60017 2128
rect 60125 2125 60175 2153
rect 60183 2125 60217 2405
rect 60341 2405 60417 2411
rect 60227 2153 60251 2377
rect 60307 2373 60331 2377
rect 60259 2169 60261 2361
rect 60263 2157 60267 2373
rect 60285 2157 60331 2373
rect 60307 2153 60331 2157
rect 60341 2153 60375 2405
rect 60125 2119 60217 2125
rect 60325 2125 60375 2153
rect 60383 2125 60417 2405
rect 60541 2405 60617 2411
rect 60427 2153 60451 2377
rect 60507 2373 60531 2377
rect 60459 2169 60461 2361
rect 60463 2157 60467 2373
rect 60485 2157 60531 2373
rect 60507 2153 60531 2157
rect 60541 2153 60575 2405
rect 60325 2119 60417 2125
rect 60525 2125 60575 2153
rect 60583 2125 60617 2405
rect 60741 2405 60817 2411
rect 60627 2153 60651 2377
rect 60707 2373 60731 2377
rect 60659 2169 60661 2361
rect 60663 2157 60667 2373
rect 60685 2157 60731 2373
rect 60707 2153 60731 2157
rect 60741 2153 60775 2405
rect 60525 2119 60617 2125
rect 60725 2125 60775 2153
rect 60783 2125 60817 2405
rect 60941 2405 61017 2411
rect 60827 2153 60851 2377
rect 60907 2373 60931 2377
rect 60859 2169 60861 2361
rect 60863 2157 60867 2373
rect 60885 2157 60931 2373
rect 60907 2153 60931 2157
rect 60941 2153 60975 2405
rect 60725 2119 60817 2125
rect 60925 2125 60975 2153
rect 60983 2125 61017 2405
rect 61027 2153 61051 2377
rect 61107 2373 61131 2377
rect 61059 2169 61061 2361
rect 61063 2157 61067 2373
rect 61085 2157 61131 2373
rect 61107 2153 61131 2157
rect 61141 2153 61417 2411
rect 61541 2411 61815 2420
rect 61943 2411 61975 2445
rect 61983 2411 62015 2445
rect 62143 2411 62175 2445
rect 62183 2411 62215 2445
rect 62343 2411 62375 2445
rect 62383 2411 62415 2445
rect 62543 2411 62575 2445
rect 62583 2411 62615 2445
rect 62743 2411 62775 2445
rect 62783 2411 62815 2445
rect 62943 2420 63215 2451
rect 63343 2461 63617 2469
rect 63343 2420 63615 2461
rect 63725 2451 63775 2479
rect 63783 2461 63817 2513
rect 63949 2479 63975 2513
rect 63783 2451 63815 2461
rect 63725 2445 63741 2451
rect 63743 2445 63815 2451
rect 63925 2451 63975 2479
rect 63983 2461 64017 2513
rect 64149 2479 64175 2513
rect 63983 2451 64015 2461
rect 63925 2445 63941 2451
rect 63943 2445 64015 2451
rect 64125 2451 64175 2479
rect 64183 2461 64217 2513
rect 64349 2479 64375 2513
rect 64183 2451 64215 2461
rect 64125 2445 64141 2451
rect 64143 2445 64215 2451
rect 64325 2451 64375 2479
rect 64383 2461 64417 2513
rect 64549 2479 64575 2513
rect 64383 2451 64415 2461
rect 64325 2445 64341 2451
rect 64343 2445 64415 2451
rect 64525 2451 64575 2479
rect 64583 2461 64617 2513
rect 64747 2479 65017 2513
rect 65147 2513 66817 2531
rect 65147 2497 65417 2513
rect 64583 2451 64615 2461
rect 64525 2445 64541 2451
rect 64543 2445 64615 2451
rect 64725 2451 65015 2479
rect 65125 2469 65417 2497
rect 65549 2479 65575 2513
rect 65125 2463 65141 2469
rect 64725 2445 64741 2451
rect 62943 2411 63217 2420
rect 61427 2162 61451 2386
rect 61507 2382 61531 2386
rect 61459 2178 61461 2370
rect 61463 2166 61467 2382
rect 61485 2166 61531 2382
rect 61507 2162 61531 2166
rect 61541 2153 61817 2411
rect 61941 2405 62017 2411
rect 61827 2153 61851 2377
rect 61907 2373 61931 2377
rect 61859 2169 61861 2361
rect 61863 2157 61867 2373
rect 61885 2157 61931 2373
rect 61907 2153 61931 2157
rect 61941 2153 61975 2405
rect 60925 2119 61017 2125
rect 61125 2128 61417 2153
rect 61525 2128 61817 2153
rect 61125 2119 61415 2128
rect 61525 2119 61541 2128
rect 61543 2119 61817 2128
rect 61925 2125 61975 2153
rect 61983 2125 62017 2405
rect 62141 2405 62217 2411
rect 62027 2153 62051 2377
rect 62107 2373 62131 2377
rect 62059 2169 62061 2361
rect 62063 2157 62067 2373
rect 62085 2157 62131 2373
rect 62107 2153 62131 2157
rect 62141 2153 62175 2405
rect 61925 2119 62017 2125
rect 62125 2125 62175 2153
rect 62183 2125 62217 2405
rect 62341 2405 62417 2411
rect 62227 2153 62251 2377
rect 62307 2373 62331 2377
rect 62259 2169 62261 2361
rect 62263 2157 62267 2373
rect 62285 2157 62331 2373
rect 62307 2153 62331 2157
rect 62341 2153 62375 2405
rect 62125 2119 62217 2125
rect 62325 2125 62375 2153
rect 62383 2125 62417 2405
rect 62541 2405 62617 2411
rect 62427 2153 62451 2377
rect 62507 2373 62531 2377
rect 62459 2169 62461 2361
rect 62463 2157 62467 2373
rect 62485 2157 62531 2373
rect 62507 2153 62531 2157
rect 62541 2153 62575 2405
rect 62325 2119 62417 2125
rect 62525 2125 62575 2153
rect 62583 2125 62617 2405
rect 62741 2405 62817 2411
rect 62627 2153 62651 2377
rect 62707 2373 62731 2377
rect 62659 2169 62661 2361
rect 62663 2157 62667 2373
rect 62685 2157 62731 2373
rect 62707 2153 62731 2157
rect 62741 2153 62775 2405
rect 62525 2119 62617 2125
rect 62725 2125 62775 2153
rect 62783 2125 62817 2405
rect 62827 2153 62851 2377
rect 62907 2373 62931 2377
rect 62859 2169 62861 2361
rect 62863 2157 62867 2373
rect 62885 2157 62931 2373
rect 62907 2153 62931 2157
rect 62941 2153 63217 2411
rect 63341 2411 63615 2420
rect 63743 2411 63775 2445
rect 63783 2411 63815 2445
rect 63943 2411 63975 2445
rect 63983 2411 64015 2445
rect 64143 2411 64175 2445
rect 64183 2411 64215 2445
rect 64343 2411 64375 2445
rect 64383 2411 64415 2445
rect 64543 2411 64575 2445
rect 64583 2411 64615 2445
rect 64743 2420 65015 2451
rect 65143 2461 65417 2469
rect 65143 2420 65415 2461
rect 65525 2451 65575 2479
rect 65583 2461 65617 2513
rect 65749 2479 65775 2513
rect 65583 2451 65615 2461
rect 65525 2445 65541 2451
rect 65543 2445 65615 2451
rect 65725 2451 65775 2479
rect 65783 2461 65817 2513
rect 65949 2479 65975 2513
rect 65783 2451 65815 2461
rect 65725 2445 65741 2451
rect 65743 2445 65815 2451
rect 65925 2451 65975 2479
rect 65983 2461 66017 2513
rect 66149 2479 66175 2513
rect 65983 2451 66015 2461
rect 65925 2445 65941 2451
rect 65943 2445 66015 2451
rect 66125 2451 66175 2479
rect 66183 2461 66217 2513
rect 66349 2479 66375 2513
rect 66183 2451 66215 2461
rect 66125 2445 66141 2451
rect 66143 2445 66215 2451
rect 66325 2451 66375 2479
rect 66383 2461 66417 2513
rect 66547 2479 66817 2513
rect 66947 2513 68617 2531
rect 66947 2497 67217 2513
rect 66383 2451 66415 2461
rect 66325 2445 66341 2451
rect 66343 2445 66415 2451
rect 66525 2451 66815 2479
rect 66925 2469 67217 2497
rect 67349 2479 67375 2513
rect 66925 2463 66941 2469
rect 66525 2445 66541 2451
rect 64743 2411 65017 2420
rect 63227 2162 63251 2386
rect 63307 2382 63331 2386
rect 63259 2178 63261 2370
rect 63263 2166 63267 2382
rect 63285 2166 63331 2382
rect 63307 2162 63331 2166
rect 63341 2153 63617 2411
rect 63741 2405 63817 2411
rect 63627 2153 63651 2377
rect 63707 2373 63731 2377
rect 63659 2169 63661 2361
rect 63663 2157 63667 2373
rect 63685 2157 63731 2373
rect 63707 2153 63731 2157
rect 63741 2153 63775 2405
rect 62725 2119 62817 2125
rect 62925 2128 63217 2153
rect 63325 2128 63617 2153
rect 62925 2119 63215 2128
rect 63325 2119 63341 2128
rect 63343 2119 63617 2128
rect 63725 2125 63775 2153
rect 63783 2125 63817 2405
rect 63941 2405 64017 2411
rect 63827 2153 63851 2377
rect 63907 2373 63931 2377
rect 63859 2169 63861 2361
rect 63863 2157 63867 2373
rect 63885 2157 63931 2373
rect 63907 2153 63931 2157
rect 63941 2153 63975 2405
rect 63725 2119 63817 2125
rect 63925 2125 63975 2153
rect 63983 2125 64017 2405
rect 64141 2405 64217 2411
rect 64027 2153 64051 2377
rect 64107 2373 64131 2377
rect 64059 2169 64061 2361
rect 64063 2157 64067 2373
rect 64085 2157 64131 2373
rect 64107 2153 64131 2157
rect 64141 2153 64175 2405
rect 63925 2119 64017 2125
rect 64125 2125 64175 2153
rect 64183 2125 64217 2405
rect 64341 2405 64417 2411
rect 64227 2153 64251 2377
rect 64307 2373 64331 2377
rect 64259 2169 64261 2361
rect 64263 2157 64267 2373
rect 64285 2157 64331 2373
rect 64307 2153 64331 2157
rect 64341 2153 64375 2405
rect 64125 2119 64217 2125
rect 64325 2125 64375 2153
rect 64383 2125 64417 2405
rect 64541 2405 64617 2411
rect 64427 2153 64451 2377
rect 64507 2373 64531 2377
rect 64459 2169 64461 2361
rect 64463 2157 64467 2373
rect 64485 2157 64531 2373
rect 64507 2153 64531 2157
rect 64541 2153 64575 2405
rect 64325 2119 64417 2125
rect 64525 2125 64575 2153
rect 64583 2125 64617 2405
rect 64627 2153 64651 2377
rect 64707 2373 64731 2377
rect 64659 2169 64661 2361
rect 64663 2157 64667 2373
rect 64685 2157 64731 2373
rect 64707 2153 64731 2157
rect 64741 2153 65017 2411
rect 65141 2411 65415 2420
rect 65543 2411 65575 2445
rect 65583 2411 65615 2445
rect 65743 2411 65775 2445
rect 65783 2411 65815 2445
rect 65943 2411 65975 2445
rect 65983 2411 66015 2445
rect 66143 2411 66175 2445
rect 66183 2411 66215 2445
rect 66343 2411 66375 2445
rect 66383 2411 66415 2445
rect 66543 2420 66815 2451
rect 66943 2461 67217 2469
rect 66943 2420 67215 2461
rect 67325 2451 67375 2479
rect 67383 2461 67417 2513
rect 67549 2479 67575 2513
rect 67383 2451 67415 2461
rect 67325 2445 67341 2451
rect 67343 2445 67415 2451
rect 67525 2451 67575 2479
rect 67583 2461 67617 2513
rect 67749 2479 67775 2513
rect 67583 2451 67615 2461
rect 67525 2445 67541 2451
rect 67543 2445 67615 2451
rect 67725 2451 67775 2479
rect 67783 2461 67817 2513
rect 67949 2479 67975 2513
rect 67783 2451 67815 2461
rect 67725 2445 67741 2451
rect 67743 2445 67815 2451
rect 67925 2451 67975 2479
rect 67983 2461 68017 2513
rect 68149 2479 68175 2513
rect 67983 2451 68015 2461
rect 67925 2445 67941 2451
rect 67943 2445 68015 2451
rect 68125 2451 68175 2479
rect 68183 2461 68217 2513
rect 68347 2479 68617 2513
rect 68183 2451 68215 2461
rect 68125 2445 68141 2451
rect 68143 2445 68215 2451
rect 68325 2451 68615 2479
rect 68725 2469 68775 2497
rect 68725 2463 68741 2469
rect 68743 2463 68811 2469
rect 68325 2445 68341 2451
rect 66543 2411 66817 2420
rect 65027 2162 65051 2386
rect 65107 2382 65131 2386
rect 65059 2178 65061 2370
rect 65063 2166 65067 2382
rect 65085 2166 65131 2382
rect 65107 2162 65131 2166
rect 65141 2153 65417 2411
rect 65541 2405 65617 2411
rect 65427 2153 65451 2377
rect 65507 2373 65531 2377
rect 65459 2169 65461 2361
rect 65463 2157 65467 2373
rect 65485 2157 65531 2373
rect 65507 2153 65531 2157
rect 65541 2153 65575 2405
rect 64525 2119 64617 2125
rect 64725 2128 65017 2153
rect 65125 2128 65417 2153
rect 64725 2119 65015 2128
rect 65125 2119 65141 2128
rect 65143 2119 65417 2128
rect 65525 2125 65575 2153
rect 65583 2125 65617 2405
rect 65741 2405 65817 2411
rect 65627 2153 65651 2377
rect 65707 2373 65731 2377
rect 65659 2169 65661 2361
rect 65663 2157 65667 2373
rect 65685 2157 65731 2373
rect 65707 2153 65731 2157
rect 65741 2153 65775 2405
rect 65525 2119 65617 2125
rect 65725 2125 65775 2153
rect 65783 2125 65817 2405
rect 65941 2405 66017 2411
rect 65827 2153 65851 2377
rect 65907 2373 65931 2377
rect 65859 2169 65861 2361
rect 65863 2157 65867 2373
rect 65885 2157 65931 2373
rect 65907 2153 65931 2157
rect 65941 2153 65975 2405
rect 65725 2119 65817 2125
rect 65925 2125 65975 2153
rect 65983 2125 66017 2405
rect 66141 2405 66217 2411
rect 66027 2153 66051 2377
rect 66107 2373 66131 2377
rect 66059 2169 66061 2361
rect 66063 2157 66067 2373
rect 66085 2157 66131 2373
rect 66107 2153 66131 2157
rect 66141 2153 66175 2405
rect 65925 2119 66017 2125
rect 66125 2125 66175 2153
rect 66183 2125 66217 2405
rect 66341 2405 66417 2411
rect 66227 2153 66251 2377
rect 66307 2373 66331 2377
rect 66259 2169 66261 2361
rect 66263 2157 66267 2373
rect 66285 2157 66331 2373
rect 66307 2153 66331 2157
rect 66341 2153 66375 2405
rect 66125 2119 66217 2125
rect 66325 2125 66375 2153
rect 66383 2125 66417 2405
rect 66427 2153 66451 2377
rect 66507 2373 66531 2377
rect 66459 2169 66461 2361
rect 66463 2157 66467 2373
rect 66485 2157 66531 2373
rect 66507 2153 66531 2157
rect 66541 2153 66817 2411
rect 66941 2411 67215 2420
rect 67343 2411 67375 2445
rect 67383 2411 67415 2445
rect 67543 2411 67575 2445
rect 67583 2411 67615 2445
rect 67743 2411 67775 2445
rect 67783 2411 67815 2445
rect 67943 2411 67975 2445
rect 67983 2411 68015 2445
rect 68143 2411 68175 2445
rect 68183 2411 68215 2445
rect 68343 2420 68615 2451
rect 68743 2429 68775 2463
rect 68799 2429 68809 2463
rect 68743 2423 68811 2429
rect 68743 2420 68775 2423
rect 68343 2411 68617 2420
rect 66827 2162 66851 2386
rect 66907 2382 66931 2386
rect 66859 2178 66861 2370
rect 66863 2166 66867 2382
rect 66885 2166 66931 2382
rect 66907 2162 66931 2166
rect 66941 2153 67217 2411
rect 67341 2405 67417 2411
rect 67227 2153 67251 2377
rect 67307 2373 67331 2377
rect 67259 2169 67261 2361
rect 67263 2157 67267 2373
rect 67285 2157 67331 2373
rect 67307 2153 67331 2157
rect 67341 2153 67375 2405
rect 66325 2119 66417 2125
rect 66525 2128 66817 2153
rect 66925 2128 67217 2153
rect 66525 2119 66815 2128
rect 66925 2119 66941 2128
rect 66943 2119 67217 2128
rect 67325 2125 67375 2153
rect 67383 2125 67417 2405
rect 67541 2405 67617 2411
rect 67427 2153 67451 2377
rect 67507 2373 67531 2377
rect 67459 2169 67461 2361
rect 67463 2157 67467 2373
rect 67485 2157 67531 2373
rect 67507 2153 67531 2157
rect 67541 2153 67575 2405
rect 67325 2119 67417 2125
rect 67525 2125 67575 2153
rect 67583 2125 67617 2405
rect 67741 2405 67817 2411
rect 67627 2153 67651 2377
rect 67707 2373 67731 2377
rect 67659 2169 67661 2361
rect 67663 2157 67667 2373
rect 67685 2157 67731 2373
rect 67707 2153 67731 2157
rect 67741 2153 67775 2405
rect 67525 2119 67617 2125
rect 67725 2125 67775 2153
rect 67783 2125 67817 2405
rect 67941 2405 68017 2411
rect 67827 2153 67851 2377
rect 67907 2373 67931 2377
rect 67859 2169 67861 2361
rect 67863 2157 67867 2373
rect 67885 2157 67931 2373
rect 67907 2153 67931 2157
rect 67941 2153 67975 2405
rect 67725 2119 67817 2125
rect 67925 2125 67975 2153
rect 67983 2125 68017 2405
rect 68141 2405 68217 2411
rect 68027 2153 68051 2377
rect 68107 2373 68131 2377
rect 68059 2169 68061 2361
rect 68063 2157 68067 2373
rect 68085 2157 68131 2373
rect 68107 2153 68131 2157
rect 68141 2153 68175 2405
rect 67925 2119 68017 2125
rect 68125 2125 68175 2153
rect 68183 2125 68217 2405
rect 68227 2153 68251 2377
rect 68307 2373 68331 2377
rect 68259 2169 68261 2361
rect 68263 2157 68267 2373
rect 68285 2157 68331 2373
rect 68307 2153 68331 2157
rect 68341 2153 68617 2411
rect 68627 2162 68651 2386
rect 68707 2382 68731 2386
rect 68659 2178 68661 2370
rect 68663 2166 68667 2382
rect 68685 2166 68731 2382
rect 68707 2162 68731 2166
rect 68741 2153 68775 2420
rect 68125 2119 68217 2125
rect 68325 2128 68617 2153
rect 68725 2128 68775 2153
rect 68325 2119 68615 2128
rect 68725 2119 68741 2128
rect 68743 2125 68775 2128
rect 68743 2119 68811 2125
rect 19943 2085 19975 2119
rect 19983 2085 20015 2119
rect 19743 2079 19815 2085
rect 19743 2069 19775 2079
rect 19183 2017 19217 2069
rect 19347 2017 19617 2069
rect 19749 2017 19775 2069
rect 19783 2069 19815 2079
rect 19943 2079 20015 2085
rect 19943 2069 19975 2079
rect 19783 2017 19817 2069
rect 19949 2017 19975 2069
rect 19983 2069 20015 2079
rect 20143 2069 20415 2119
rect 20543 2085 20575 2119
rect 20583 2085 20615 2119
rect 20543 2079 20615 2085
rect 20543 2069 20575 2079
rect 19983 2017 20017 2069
rect 20147 2017 20417 2069
rect 20549 2017 20575 2069
rect 20583 2069 20615 2079
rect 20743 2085 20775 2119
rect 20783 2085 20815 2119
rect 20743 2079 20815 2085
rect 20743 2069 20775 2079
rect 20583 2017 20617 2069
rect 20749 2017 20775 2069
rect 20783 2069 20815 2079
rect 20943 2085 20975 2119
rect 20983 2085 21015 2119
rect 20943 2079 21015 2085
rect 20943 2069 20975 2079
rect 20783 2017 20817 2069
rect 20949 2017 20975 2069
rect 20983 2069 21015 2079
rect 21143 2085 21175 2119
rect 21183 2085 21215 2119
rect 21143 2079 21215 2085
rect 21143 2069 21175 2079
rect 20983 2017 21017 2069
rect 21149 2017 21175 2069
rect 21183 2069 21215 2079
rect 21343 2085 21375 2119
rect 21383 2085 21415 2119
rect 21343 2079 21415 2085
rect 21343 2069 21375 2079
rect 21183 2017 21217 2069
rect 21349 2017 21375 2069
rect 21383 2069 21415 2079
rect 21543 2069 21815 2119
rect 21943 2069 22215 2119
rect 22343 2085 22375 2119
rect 22383 2085 22415 2119
rect 22343 2079 22415 2085
rect 22343 2069 22375 2079
rect 21383 2017 21417 2069
rect 21547 2017 21817 2069
rect 21947 2017 22217 2069
rect 22349 2017 22375 2069
rect 22383 2069 22415 2079
rect 22543 2085 22575 2119
rect 22583 2085 22615 2119
rect 22543 2079 22615 2085
rect 22543 2069 22575 2079
rect 22383 2017 22417 2069
rect 22549 2017 22575 2069
rect 22583 2069 22615 2079
rect 22743 2085 22775 2119
rect 22783 2085 22815 2119
rect 22743 2079 22815 2085
rect 22743 2069 22775 2079
rect 22583 2017 22617 2069
rect 22749 2017 22775 2069
rect 22783 2069 22815 2079
rect 22943 2085 22975 2119
rect 22983 2085 23015 2119
rect 22943 2079 23015 2085
rect 22943 2069 22975 2079
rect 22783 2017 22817 2069
rect 22949 2017 22975 2069
rect 22983 2069 23015 2079
rect 23143 2085 23175 2119
rect 23183 2085 23215 2119
rect 23143 2079 23215 2085
rect 23143 2069 23175 2079
rect 22983 2017 23017 2069
rect 23149 2017 23175 2069
rect 23183 2069 23215 2079
rect 23343 2069 23615 2119
rect 23743 2069 24015 2119
rect 24143 2085 24175 2119
rect 24183 2085 24215 2119
rect 24143 2079 24215 2085
rect 24143 2069 24175 2079
rect 23183 2017 23217 2069
rect 23347 2017 23617 2069
rect 23747 2017 24017 2069
rect 24149 2017 24175 2069
rect 24183 2069 24215 2079
rect 24343 2085 24375 2119
rect 24383 2085 24415 2119
rect 24343 2079 24415 2085
rect 24343 2069 24375 2079
rect 24183 2017 24217 2069
rect 24349 2017 24375 2069
rect 24383 2069 24415 2079
rect 24543 2085 24575 2119
rect 24583 2085 24615 2119
rect 24543 2079 24615 2085
rect 24543 2069 24575 2079
rect 24383 2017 24417 2069
rect 24549 2017 24575 2069
rect 24583 2069 24615 2079
rect 24743 2085 24775 2119
rect 24783 2085 24815 2119
rect 24743 2079 24815 2085
rect 24743 2069 24775 2079
rect 24583 2017 24617 2069
rect 24749 2017 24775 2069
rect 24783 2069 24815 2079
rect 24943 2085 24975 2119
rect 24983 2085 25015 2119
rect 24943 2079 25015 2085
rect 24943 2069 24975 2079
rect 24783 2017 24817 2069
rect 24949 2017 24975 2069
rect 24983 2069 25015 2079
rect 25143 2069 25415 2119
rect 25543 2069 25815 2119
rect 25943 2085 25975 2119
rect 25983 2085 26015 2119
rect 25943 2079 26015 2085
rect 25943 2069 25975 2079
rect 24983 2017 25017 2069
rect 25147 2017 25417 2069
rect 25547 2017 25817 2069
rect 25949 2017 25975 2069
rect 25983 2069 26015 2079
rect 26143 2085 26175 2119
rect 26183 2085 26215 2119
rect 26143 2079 26215 2085
rect 26143 2069 26175 2079
rect 25983 2017 26017 2069
rect 26149 2017 26175 2069
rect 26183 2069 26215 2079
rect 26343 2085 26375 2119
rect 26383 2085 26415 2119
rect 26343 2079 26415 2085
rect 26343 2069 26375 2079
rect 26183 2017 26217 2069
rect 26349 2017 26375 2069
rect 26383 2069 26415 2079
rect 26543 2085 26575 2119
rect 26583 2085 26615 2119
rect 26543 2079 26615 2085
rect 26543 2069 26575 2079
rect 26383 2017 26417 2069
rect 26549 2017 26575 2069
rect 26583 2069 26615 2079
rect 26743 2085 26775 2119
rect 26783 2085 26815 2119
rect 26743 2079 26815 2085
rect 26743 2069 26775 2079
rect 26583 2017 26617 2069
rect 26749 2017 26775 2069
rect 26783 2069 26815 2079
rect 26943 2069 27215 2119
rect 27343 2069 27615 2119
rect 27743 2085 27775 2119
rect 27783 2085 27815 2119
rect 27743 2079 27815 2085
rect 27743 2069 27775 2079
rect 26783 2017 26817 2069
rect 26947 2017 27217 2069
rect 27347 2017 27617 2069
rect 27749 2017 27775 2069
rect 27783 2069 27815 2079
rect 27943 2085 27975 2119
rect 27983 2085 28015 2119
rect 27943 2079 28015 2085
rect 27943 2069 27975 2079
rect 27783 2017 27817 2069
rect 27949 2017 27975 2069
rect 27983 2069 28015 2079
rect 28143 2085 28175 2119
rect 28183 2085 28215 2119
rect 28143 2079 28215 2085
rect 28143 2069 28175 2079
rect 27983 2017 28017 2069
rect 28149 2017 28175 2069
rect 28183 2069 28215 2079
rect 28343 2085 28375 2119
rect 28383 2085 28415 2119
rect 28343 2079 28415 2085
rect 28343 2069 28375 2079
rect 28183 2017 28217 2069
rect 28349 2017 28375 2069
rect 28383 2069 28415 2079
rect 28543 2085 28575 2119
rect 28583 2085 28615 2119
rect 28543 2079 28615 2085
rect 28543 2069 28575 2079
rect 28383 2017 28417 2069
rect 28549 2017 28575 2069
rect 28583 2069 28615 2079
rect 28743 2069 29015 2119
rect 29143 2069 29415 2119
rect 29543 2085 29575 2119
rect 29583 2085 29615 2119
rect 29543 2079 29615 2085
rect 29543 2069 29575 2079
rect 28583 2017 28617 2069
rect 28747 2017 29017 2069
rect 29147 2017 29417 2069
rect 29549 2017 29575 2069
rect 29583 2069 29615 2079
rect 29743 2085 29775 2119
rect 29783 2085 29815 2119
rect 29743 2079 29815 2085
rect 29743 2069 29775 2079
rect 29583 2017 29617 2069
rect 29749 2017 29775 2069
rect 29783 2069 29815 2079
rect 29943 2085 29975 2119
rect 29983 2085 30015 2119
rect 29943 2079 30015 2085
rect 29943 2069 29975 2079
rect 29783 2017 29817 2069
rect 29949 2017 29975 2069
rect 29983 2069 30015 2079
rect 30143 2085 30175 2119
rect 30183 2085 30215 2119
rect 30143 2079 30215 2085
rect 30143 2069 30175 2079
rect 29983 2017 30017 2069
rect 30149 2017 30175 2069
rect 30183 2069 30215 2079
rect 30343 2085 30375 2119
rect 30383 2085 30415 2119
rect 30343 2079 30415 2085
rect 30343 2069 30375 2079
rect 30183 2017 30217 2069
rect 30349 2017 30375 2069
rect 30383 2069 30415 2079
rect 30543 2069 30815 2119
rect 30943 2069 31215 2119
rect 31343 2085 31375 2119
rect 31383 2085 31415 2119
rect 31343 2079 31415 2085
rect 31343 2069 31375 2079
rect 30383 2017 30417 2069
rect 30547 2017 30817 2069
rect 30947 2017 31217 2069
rect 31349 2017 31375 2069
rect 31383 2069 31415 2079
rect 31543 2085 31575 2119
rect 31583 2085 31615 2119
rect 31543 2079 31615 2085
rect 31543 2069 31575 2079
rect 31383 2017 31417 2069
rect 31549 2017 31575 2069
rect 31583 2069 31615 2079
rect 31743 2085 31775 2119
rect 31783 2085 31815 2119
rect 31743 2079 31815 2085
rect 31743 2069 31775 2079
rect 31583 2017 31617 2069
rect 31749 2017 31775 2069
rect 31783 2069 31815 2079
rect 31943 2085 31975 2119
rect 31983 2085 32015 2119
rect 31943 2079 32015 2085
rect 31943 2069 31975 2079
rect 31783 2017 31817 2069
rect 31949 2017 31975 2069
rect 31983 2069 32015 2079
rect 32143 2085 32175 2119
rect 32183 2085 32215 2119
rect 32143 2079 32215 2085
rect 32143 2069 32175 2079
rect 31983 2017 32017 2069
rect 32149 2017 32175 2069
rect 32183 2069 32215 2079
rect 32343 2069 32615 2119
rect 32743 2069 33015 2119
rect 33143 2085 33175 2119
rect 33183 2085 33215 2119
rect 33143 2079 33215 2085
rect 33143 2069 33175 2079
rect 32183 2017 32217 2069
rect 32347 2017 32617 2069
rect 32747 2017 33017 2069
rect 33149 2017 33175 2069
rect 33183 2069 33215 2079
rect 33343 2085 33375 2119
rect 33383 2085 33415 2119
rect 33343 2079 33415 2085
rect 33343 2069 33375 2079
rect 33183 2017 33217 2069
rect 33349 2017 33375 2069
rect 33383 2069 33415 2079
rect 33543 2085 33575 2119
rect 33583 2085 33615 2119
rect 33543 2079 33615 2085
rect 33543 2069 33575 2079
rect 33383 2017 33417 2069
rect 33549 2017 33575 2069
rect 33583 2069 33615 2079
rect 33743 2085 33775 2119
rect 33783 2085 33815 2119
rect 33743 2079 33815 2085
rect 33743 2069 33775 2079
rect 33583 2017 33617 2069
rect 33749 2017 33775 2069
rect 33783 2069 33815 2079
rect 33943 2085 33975 2119
rect 33983 2085 34015 2119
rect 33943 2079 34015 2085
rect 33943 2069 33975 2079
rect 33783 2017 33817 2069
rect 33949 2017 33975 2069
rect 33983 2069 34015 2079
rect 34143 2069 34415 2119
rect 34543 2069 34815 2119
rect 34943 2085 34975 2119
rect 34983 2085 35015 2119
rect 34943 2079 35015 2085
rect 34943 2069 34975 2079
rect 33983 2017 34017 2069
rect 34147 2017 34417 2069
rect 34547 2017 34817 2069
rect 34949 2017 34975 2069
rect 34983 2069 35015 2079
rect 35143 2085 35175 2119
rect 35183 2085 35215 2119
rect 35143 2079 35215 2085
rect 35143 2069 35175 2079
rect 34983 2017 35017 2069
rect 35149 2017 35175 2069
rect 35183 2069 35215 2079
rect 35343 2085 35375 2119
rect 35383 2085 35415 2119
rect 35343 2079 35415 2085
rect 35343 2069 35375 2079
rect 35183 2017 35217 2069
rect 35349 2017 35375 2069
rect 35383 2069 35415 2079
rect 35543 2085 35575 2119
rect 35583 2085 35615 2119
rect 35543 2079 35615 2085
rect 35543 2069 35575 2079
rect 35383 2017 35417 2069
rect 35549 2017 35575 2069
rect 35583 2069 35615 2079
rect 35743 2085 35775 2119
rect 35783 2085 35815 2119
rect 35743 2079 35815 2085
rect 35743 2069 35775 2079
rect 35583 2017 35617 2069
rect 35749 2017 35775 2069
rect 35783 2069 35815 2079
rect 35943 2069 36215 2119
rect 36343 2069 36615 2119
rect 36743 2085 36775 2119
rect 36783 2085 36815 2119
rect 36743 2079 36815 2085
rect 36743 2069 36775 2079
rect 35783 2017 35817 2069
rect 35947 2017 36217 2069
rect 36347 2017 36617 2069
rect 36749 2017 36775 2069
rect 36783 2069 36815 2079
rect 36943 2085 36975 2119
rect 36983 2085 37015 2119
rect 36943 2079 37015 2085
rect 36943 2069 36975 2079
rect 36783 2017 36817 2069
rect 36949 2017 36975 2069
rect 36983 2069 37015 2079
rect 37143 2085 37175 2119
rect 37183 2085 37215 2119
rect 37143 2079 37215 2085
rect 37143 2069 37175 2079
rect 36983 2017 37017 2069
rect 37149 2017 37175 2069
rect 37183 2069 37215 2079
rect 37343 2085 37375 2119
rect 37383 2085 37415 2119
rect 37343 2079 37415 2085
rect 37343 2069 37375 2079
rect 37183 2017 37217 2069
rect 37349 2017 37375 2069
rect 37383 2069 37415 2079
rect 37543 2085 37575 2119
rect 37583 2085 37615 2119
rect 37543 2079 37615 2085
rect 37543 2069 37575 2079
rect 37383 2017 37417 2069
rect 37549 2017 37575 2069
rect 37583 2069 37615 2079
rect 37743 2069 38015 2119
rect 38143 2069 38415 2119
rect 38543 2085 38575 2119
rect 38583 2085 38615 2119
rect 38543 2079 38615 2085
rect 38543 2069 38575 2079
rect 37583 2017 37617 2069
rect 37747 2017 38017 2069
rect 38147 2017 38417 2069
rect 38549 2017 38575 2069
rect 38583 2069 38615 2079
rect 38743 2085 38775 2119
rect 38783 2085 38815 2119
rect 38743 2079 38815 2085
rect 38743 2069 38775 2079
rect 38583 2017 38617 2069
rect 38749 2017 38775 2069
rect 38783 2069 38815 2079
rect 38943 2085 38975 2119
rect 38983 2085 39015 2119
rect 38943 2079 39015 2085
rect 38943 2069 38975 2079
rect 38783 2017 38817 2069
rect 38949 2017 38975 2069
rect 38983 2069 39015 2079
rect 39143 2085 39175 2119
rect 39183 2085 39215 2119
rect 39143 2079 39215 2085
rect 39143 2069 39175 2079
rect 38983 2017 39017 2069
rect 39149 2017 39175 2069
rect 39183 2069 39215 2079
rect 39343 2085 39375 2119
rect 39383 2085 39415 2119
rect 39343 2079 39415 2085
rect 39343 2069 39375 2079
rect 39183 2017 39217 2069
rect 39349 2017 39375 2069
rect 39383 2069 39415 2079
rect 39543 2069 39815 2119
rect 39943 2069 40215 2119
rect 40343 2085 40375 2119
rect 40383 2085 40415 2119
rect 40343 2079 40415 2085
rect 40343 2069 40375 2079
rect 39383 2017 39417 2069
rect 39547 2017 39817 2069
rect 39947 2017 40217 2069
rect 40349 2017 40375 2069
rect 40383 2069 40415 2079
rect 40543 2085 40575 2119
rect 40583 2085 40615 2119
rect 40543 2079 40615 2085
rect 40543 2069 40575 2079
rect 40383 2017 40417 2069
rect 40549 2017 40575 2069
rect 40583 2069 40615 2079
rect 40743 2085 40775 2119
rect 40783 2085 40815 2119
rect 40743 2079 40815 2085
rect 40743 2069 40775 2079
rect 40583 2017 40617 2069
rect 40749 2017 40775 2069
rect 40783 2069 40815 2079
rect 40943 2085 40975 2119
rect 40983 2085 41015 2119
rect 40943 2079 41015 2085
rect 40943 2069 40975 2079
rect 40783 2017 40817 2069
rect 40949 2017 40975 2069
rect 40983 2069 41015 2079
rect 41143 2085 41175 2119
rect 41183 2085 41215 2119
rect 41143 2079 41215 2085
rect 41143 2069 41175 2079
rect 40983 2017 41017 2069
rect 41149 2017 41175 2069
rect 41183 2069 41215 2079
rect 41343 2069 41615 2119
rect 41743 2069 42015 2119
rect 42143 2085 42175 2119
rect 42183 2085 42215 2119
rect 42143 2079 42215 2085
rect 42143 2069 42175 2079
rect 41183 2017 41217 2069
rect 41347 2017 41617 2069
rect 41747 2017 42017 2069
rect 42149 2017 42175 2069
rect 42183 2069 42215 2079
rect 42343 2085 42375 2119
rect 42383 2085 42415 2119
rect 42343 2079 42415 2085
rect 42343 2069 42375 2079
rect 42183 2017 42217 2069
rect 42349 2017 42375 2069
rect 42383 2069 42415 2079
rect 42543 2085 42575 2119
rect 42583 2085 42615 2119
rect 42543 2079 42615 2085
rect 42543 2069 42575 2079
rect 42383 2017 42417 2069
rect 42549 2017 42575 2069
rect 42583 2069 42615 2079
rect 42743 2085 42775 2119
rect 42783 2085 42815 2119
rect 42743 2079 42815 2085
rect 42743 2069 42775 2079
rect 42583 2017 42617 2069
rect 42749 2017 42775 2069
rect 42783 2069 42815 2079
rect 42943 2085 42975 2119
rect 42983 2085 43015 2119
rect 42943 2079 43015 2085
rect 42943 2069 42975 2079
rect 42783 2017 42817 2069
rect 42949 2017 42975 2069
rect 42983 2069 43015 2079
rect 43143 2069 43415 2119
rect 43543 2069 43815 2119
rect 43943 2085 43975 2119
rect 43983 2085 44015 2119
rect 43943 2079 44015 2085
rect 43943 2069 43975 2079
rect 42983 2017 43017 2069
rect 43147 2017 43417 2069
rect 43547 2017 43817 2069
rect 43949 2017 43975 2069
rect 43983 2069 44015 2079
rect 44143 2085 44175 2119
rect 44183 2085 44215 2119
rect 44143 2079 44215 2085
rect 44143 2069 44175 2079
rect 43983 2017 44017 2069
rect 44149 2017 44175 2069
rect 44183 2069 44215 2079
rect 44343 2085 44375 2119
rect 44383 2085 44415 2119
rect 44343 2079 44415 2085
rect 44343 2069 44375 2079
rect 44183 2017 44217 2069
rect 44349 2017 44375 2069
rect 44383 2069 44415 2079
rect 44543 2085 44575 2119
rect 44583 2085 44615 2119
rect 44543 2079 44615 2085
rect 44543 2069 44575 2079
rect 44383 2017 44417 2069
rect 44549 2017 44575 2069
rect 44583 2069 44615 2079
rect 44743 2085 44775 2119
rect 44783 2085 44815 2119
rect 44743 2079 44815 2085
rect 44743 2069 44775 2079
rect 44583 2017 44617 2069
rect 44749 2017 44775 2069
rect 44783 2069 44815 2079
rect 44943 2069 45215 2119
rect 45343 2069 45615 2119
rect 45743 2085 45775 2119
rect 45783 2085 45815 2119
rect 45743 2079 45815 2085
rect 45743 2069 45775 2079
rect 44783 2017 44817 2069
rect 44947 2017 45217 2069
rect 45347 2017 45617 2069
rect 45749 2017 45775 2069
rect 45783 2069 45815 2079
rect 45943 2085 45975 2119
rect 45983 2085 46015 2119
rect 45943 2079 46015 2085
rect 45943 2069 45975 2079
rect 45783 2017 45817 2069
rect 45949 2017 45975 2069
rect 45983 2069 46015 2079
rect 46143 2085 46175 2119
rect 46183 2085 46215 2119
rect 46143 2079 46215 2085
rect 46143 2069 46175 2079
rect 45983 2017 46017 2069
rect 46149 2017 46175 2069
rect 46183 2069 46215 2079
rect 46343 2085 46375 2119
rect 46383 2085 46415 2119
rect 46343 2079 46415 2085
rect 46343 2069 46375 2079
rect 46183 2017 46217 2069
rect 46349 2017 46375 2069
rect 46383 2069 46415 2079
rect 46543 2085 46575 2119
rect 46583 2085 46615 2119
rect 46543 2079 46615 2085
rect 46543 2069 46575 2079
rect 46383 2017 46417 2069
rect 46549 2017 46575 2069
rect 46583 2069 46615 2079
rect 46743 2069 47015 2119
rect 47143 2069 47415 2119
rect 47543 2085 47575 2119
rect 47583 2085 47615 2119
rect 47543 2079 47615 2085
rect 47543 2069 47575 2079
rect 46583 2017 46617 2069
rect 46747 2017 47017 2069
rect 47147 2017 47417 2069
rect 47549 2017 47575 2069
rect 47583 2069 47615 2079
rect 47743 2085 47775 2119
rect 47783 2085 47815 2119
rect 47743 2079 47815 2085
rect 47743 2069 47775 2079
rect 47583 2017 47617 2069
rect 47749 2017 47775 2069
rect 47783 2069 47815 2079
rect 47943 2085 47975 2119
rect 47983 2085 48015 2119
rect 47943 2079 48015 2085
rect 47943 2069 47975 2079
rect 47783 2017 47817 2069
rect 47949 2017 47975 2069
rect 47983 2069 48015 2079
rect 48143 2085 48175 2119
rect 48183 2085 48215 2119
rect 48143 2079 48215 2085
rect 48143 2069 48175 2079
rect 47983 2017 48017 2069
rect 48149 2017 48175 2069
rect 48183 2069 48215 2079
rect 48343 2085 48375 2119
rect 48383 2085 48415 2119
rect 48343 2079 48415 2085
rect 48343 2069 48375 2079
rect 48183 2017 48217 2069
rect 48349 2017 48375 2069
rect 48383 2069 48415 2079
rect 48543 2069 48815 2119
rect 48943 2069 49215 2119
rect 49343 2085 49375 2119
rect 49383 2085 49415 2119
rect 49343 2079 49415 2085
rect 49343 2069 49375 2079
rect 48383 2017 48417 2069
rect 48547 2017 48817 2069
rect 48947 2017 49217 2069
rect 49349 2017 49375 2069
rect 49383 2069 49415 2079
rect 49543 2085 49575 2119
rect 49583 2085 49615 2119
rect 49543 2079 49615 2085
rect 49543 2069 49575 2079
rect 49383 2017 49417 2069
rect 49549 2017 49575 2069
rect 49583 2069 49615 2079
rect 49743 2085 49775 2119
rect 49783 2085 49815 2119
rect 49743 2079 49815 2085
rect 49743 2069 49775 2079
rect 49583 2017 49617 2069
rect 49749 2017 49775 2069
rect 49783 2069 49815 2079
rect 49943 2085 49975 2119
rect 49983 2085 50015 2119
rect 49943 2079 50015 2085
rect 49943 2069 49975 2079
rect 49783 2017 49817 2069
rect 49949 2017 49975 2069
rect 49983 2069 50015 2079
rect 50143 2085 50175 2119
rect 50183 2085 50215 2119
rect 50143 2079 50215 2085
rect 50143 2069 50175 2079
rect 49983 2017 50017 2069
rect 50149 2017 50175 2069
rect 50183 2069 50215 2079
rect 50343 2069 50615 2119
rect 50743 2069 51015 2119
rect 51143 2085 51175 2119
rect 51183 2085 51215 2119
rect 51143 2079 51215 2085
rect 51143 2069 51175 2079
rect 50183 2017 50217 2069
rect 50347 2017 50617 2069
rect 50747 2017 51017 2069
rect 51149 2017 51175 2069
rect 51183 2069 51215 2079
rect 51343 2085 51375 2119
rect 51383 2085 51415 2119
rect 51343 2079 51415 2085
rect 51343 2069 51375 2079
rect 51183 2017 51217 2069
rect 51349 2017 51375 2069
rect 51383 2069 51415 2079
rect 51543 2085 51575 2119
rect 51583 2085 51615 2119
rect 51543 2079 51615 2085
rect 51543 2069 51575 2079
rect 51383 2017 51417 2069
rect 51549 2017 51575 2069
rect 51583 2069 51615 2079
rect 51743 2085 51775 2119
rect 51783 2085 51815 2119
rect 51743 2079 51815 2085
rect 51743 2069 51775 2079
rect 51583 2017 51617 2069
rect 51749 2017 51775 2069
rect 51783 2069 51815 2079
rect 51943 2085 51975 2119
rect 51983 2085 52015 2119
rect 51943 2079 52015 2085
rect 51943 2069 51975 2079
rect 51783 2017 51817 2069
rect 51949 2017 51975 2069
rect 51983 2069 52015 2079
rect 52143 2069 52415 2119
rect 52543 2069 52815 2119
rect 52943 2085 52975 2119
rect 52983 2085 53015 2119
rect 52943 2079 53015 2085
rect 52943 2069 52975 2079
rect 51983 2017 52017 2069
rect 52147 2017 52417 2069
rect 52547 2017 52817 2069
rect 52949 2017 52975 2069
rect 52983 2069 53015 2079
rect 53143 2085 53175 2119
rect 53183 2085 53215 2119
rect 53143 2079 53215 2085
rect 53143 2069 53175 2079
rect 52983 2017 53017 2069
rect 53149 2017 53175 2069
rect 53183 2069 53215 2079
rect 53343 2085 53375 2119
rect 53383 2085 53415 2119
rect 53343 2079 53415 2085
rect 53343 2069 53375 2079
rect 53183 2017 53217 2069
rect 53349 2017 53375 2069
rect 53383 2069 53415 2079
rect 53543 2085 53575 2119
rect 53583 2085 53615 2119
rect 53543 2079 53615 2085
rect 53543 2069 53575 2079
rect 53383 2017 53417 2069
rect 53549 2017 53575 2069
rect 53583 2069 53615 2079
rect 53743 2085 53775 2119
rect 53783 2085 53815 2119
rect 53743 2079 53815 2085
rect 53743 2069 53775 2079
rect 53583 2017 53617 2069
rect 53749 2017 53775 2069
rect 53783 2069 53815 2079
rect 53943 2069 54215 2119
rect 54343 2069 54615 2119
rect 54743 2085 54775 2119
rect 54783 2085 54815 2119
rect 54743 2079 54815 2085
rect 54743 2069 54775 2079
rect 53783 2017 53817 2069
rect 53947 2017 54217 2069
rect 54347 2017 54617 2069
rect 54749 2017 54775 2069
rect 54783 2069 54815 2079
rect 54943 2085 54975 2119
rect 54983 2085 55015 2119
rect 54943 2079 55015 2085
rect 54943 2069 54975 2079
rect 54783 2017 54817 2069
rect 54949 2017 54975 2069
rect 54983 2069 55015 2079
rect 55143 2085 55175 2119
rect 55183 2085 55215 2119
rect 55143 2079 55215 2085
rect 55143 2069 55175 2079
rect 54983 2017 55017 2069
rect 55149 2017 55175 2069
rect 55183 2069 55215 2079
rect 55343 2085 55375 2119
rect 55383 2085 55415 2119
rect 55343 2079 55415 2085
rect 55343 2069 55375 2079
rect 55183 2017 55217 2069
rect 55349 2017 55375 2069
rect 55383 2069 55415 2079
rect 55543 2085 55575 2119
rect 55583 2085 55615 2119
rect 55543 2079 55615 2085
rect 55543 2069 55575 2079
rect 55383 2017 55417 2069
rect 55549 2017 55575 2069
rect 55583 2069 55615 2079
rect 55743 2069 56015 2119
rect 56143 2069 56415 2119
rect 56543 2085 56575 2119
rect 56583 2085 56615 2119
rect 56543 2079 56615 2085
rect 56543 2069 56575 2079
rect 55583 2017 55617 2069
rect 55747 2017 56017 2069
rect 56147 2017 56417 2069
rect 56549 2017 56575 2069
rect 56583 2069 56615 2079
rect 56743 2085 56775 2119
rect 56783 2085 56815 2119
rect 56743 2079 56815 2085
rect 56743 2069 56775 2079
rect 56583 2017 56617 2069
rect 56749 2017 56775 2069
rect 56783 2069 56815 2079
rect 56943 2085 56975 2119
rect 56983 2085 57015 2119
rect 56943 2079 57015 2085
rect 56943 2069 56975 2079
rect 56783 2017 56817 2069
rect 56949 2017 56975 2069
rect 56983 2069 57015 2079
rect 57143 2085 57175 2119
rect 57183 2085 57215 2119
rect 57143 2079 57215 2085
rect 57143 2069 57175 2079
rect 56983 2017 57017 2069
rect 57149 2017 57175 2069
rect 57183 2069 57215 2079
rect 57343 2085 57375 2119
rect 57383 2085 57415 2119
rect 57343 2079 57415 2085
rect 57343 2069 57375 2079
rect 57183 2017 57217 2069
rect 57349 2017 57375 2069
rect 57383 2069 57415 2079
rect 57543 2069 57815 2119
rect 57943 2069 58215 2119
rect 58343 2085 58375 2119
rect 58383 2085 58415 2119
rect 58343 2079 58415 2085
rect 58343 2069 58375 2079
rect 57383 2017 57417 2069
rect 57547 2017 57817 2069
rect 57947 2017 58217 2069
rect 58349 2017 58375 2069
rect 58383 2069 58415 2079
rect 58543 2085 58575 2119
rect 58583 2085 58615 2119
rect 58543 2079 58615 2085
rect 58543 2069 58575 2079
rect 58383 2017 58417 2069
rect 58549 2017 58575 2069
rect 58583 2069 58615 2079
rect 58743 2085 58775 2119
rect 58783 2085 58815 2119
rect 58743 2079 58815 2085
rect 58743 2069 58775 2079
rect 58583 2017 58617 2069
rect 58749 2017 58775 2069
rect 58783 2069 58815 2079
rect 58943 2085 58975 2119
rect 58983 2085 59015 2119
rect 58943 2079 59015 2085
rect 58943 2069 58975 2079
rect 58783 2017 58817 2069
rect 58949 2017 58975 2069
rect 58983 2069 59015 2079
rect 59143 2085 59175 2119
rect 59183 2085 59215 2119
rect 59143 2079 59215 2085
rect 59143 2069 59175 2079
rect 58983 2017 59017 2069
rect 59149 2017 59175 2069
rect 59183 2069 59215 2079
rect 59343 2069 59615 2119
rect 59743 2069 60015 2119
rect 60143 2085 60175 2119
rect 60183 2085 60215 2119
rect 60143 2079 60215 2085
rect 60143 2069 60175 2079
rect 59183 2017 59217 2069
rect 59347 2017 59617 2069
rect 59747 2017 60017 2069
rect 60149 2017 60175 2069
rect 60183 2069 60215 2079
rect 60343 2085 60375 2119
rect 60383 2085 60415 2119
rect 60343 2079 60415 2085
rect 60343 2069 60375 2079
rect 60183 2017 60217 2069
rect 60349 2017 60375 2069
rect 60383 2069 60415 2079
rect 60543 2085 60575 2119
rect 60583 2085 60615 2119
rect 60543 2079 60615 2085
rect 60543 2069 60575 2079
rect 60383 2017 60417 2069
rect 60549 2017 60575 2069
rect 60583 2069 60615 2079
rect 60743 2085 60775 2119
rect 60783 2085 60815 2119
rect 60743 2079 60815 2085
rect 60743 2069 60775 2079
rect 60583 2017 60617 2069
rect 60749 2017 60775 2069
rect 60783 2069 60815 2079
rect 60943 2085 60975 2119
rect 60983 2085 61015 2119
rect 60943 2079 61015 2085
rect 60943 2069 60975 2079
rect 60783 2017 60817 2069
rect 60949 2017 60975 2069
rect 60983 2069 61015 2079
rect 61143 2069 61415 2119
rect 61543 2069 61815 2119
rect 61943 2085 61975 2119
rect 61983 2085 62015 2119
rect 61943 2079 62015 2085
rect 61943 2069 61975 2079
rect 60983 2017 61017 2069
rect 61147 2017 61417 2069
rect 61547 2017 61817 2069
rect 61949 2017 61975 2069
rect 61983 2069 62015 2079
rect 62143 2085 62175 2119
rect 62183 2085 62215 2119
rect 62143 2079 62215 2085
rect 62143 2069 62175 2079
rect 61983 2017 62017 2069
rect 62149 2017 62175 2069
rect 62183 2069 62215 2079
rect 62343 2085 62375 2119
rect 62383 2085 62415 2119
rect 62343 2079 62415 2085
rect 62343 2069 62375 2079
rect 62183 2017 62217 2069
rect 62349 2017 62375 2069
rect 62383 2069 62415 2079
rect 62543 2085 62575 2119
rect 62583 2085 62615 2119
rect 62543 2079 62615 2085
rect 62543 2069 62575 2079
rect 62383 2017 62417 2069
rect 62549 2017 62575 2069
rect 62583 2069 62615 2079
rect 62743 2085 62775 2119
rect 62783 2085 62815 2119
rect 62743 2079 62815 2085
rect 62743 2069 62775 2079
rect 62583 2017 62617 2069
rect 62749 2017 62775 2069
rect 62783 2069 62815 2079
rect 62943 2069 63215 2119
rect 63343 2069 63615 2119
rect 63743 2085 63775 2119
rect 63783 2085 63815 2119
rect 63743 2079 63815 2085
rect 63743 2069 63775 2079
rect 62783 2017 62817 2069
rect 62947 2017 63217 2069
rect 63347 2017 63617 2069
rect 63749 2017 63775 2069
rect 63783 2069 63815 2079
rect 63943 2085 63975 2119
rect 63983 2085 64015 2119
rect 63943 2079 64015 2085
rect 63943 2069 63975 2079
rect 63783 2017 63817 2069
rect 63949 2017 63975 2069
rect 63983 2069 64015 2079
rect 64143 2085 64175 2119
rect 64183 2085 64215 2119
rect 64143 2079 64215 2085
rect 64143 2069 64175 2079
rect 63983 2017 64017 2069
rect 64149 2017 64175 2069
rect 64183 2069 64215 2079
rect 64343 2085 64375 2119
rect 64383 2085 64415 2119
rect 64343 2079 64415 2085
rect 64343 2069 64375 2079
rect 64183 2017 64217 2069
rect 64349 2017 64375 2069
rect 64383 2069 64415 2079
rect 64543 2085 64575 2119
rect 64583 2085 64615 2119
rect 64543 2079 64615 2085
rect 64543 2069 64575 2079
rect 64383 2017 64417 2069
rect 64549 2017 64575 2069
rect 64583 2069 64615 2079
rect 64743 2069 65015 2119
rect 65143 2069 65415 2119
rect 65543 2085 65575 2119
rect 65583 2085 65615 2119
rect 65543 2079 65615 2085
rect 65543 2069 65575 2079
rect 64583 2017 64617 2069
rect 64747 2017 65017 2069
rect 65147 2017 65417 2069
rect 65549 2017 65575 2069
rect 65583 2069 65615 2079
rect 65743 2085 65775 2119
rect 65783 2085 65815 2119
rect 65743 2079 65815 2085
rect 65743 2069 65775 2079
rect 65583 2017 65617 2069
rect 65749 2017 65775 2069
rect 65783 2069 65815 2079
rect 65943 2085 65975 2119
rect 65983 2085 66015 2119
rect 65943 2079 66015 2085
rect 65943 2069 65975 2079
rect 65783 2017 65817 2069
rect 65949 2017 65975 2069
rect 65983 2069 66015 2079
rect 66143 2085 66175 2119
rect 66183 2085 66215 2119
rect 66143 2079 66215 2085
rect 66143 2069 66175 2079
rect 65983 2017 66017 2069
rect 66149 2017 66175 2069
rect 66183 2069 66215 2079
rect 66343 2085 66375 2119
rect 66383 2085 66415 2119
rect 66343 2079 66415 2085
rect 66343 2069 66375 2079
rect 66183 2017 66217 2069
rect 66349 2017 66375 2069
rect 66383 2069 66415 2079
rect 66543 2069 66815 2119
rect 66943 2069 67215 2119
rect 67343 2085 67375 2119
rect 67383 2085 67415 2119
rect 67343 2079 67415 2085
rect 67343 2069 67375 2079
rect 66383 2017 66417 2069
rect 66547 2017 66817 2069
rect 66947 2017 67217 2069
rect 67349 2017 67375 2069
rect 67383 2069 67415 2079
rect 67543 2085 67575 2119
rect 67583 2085 67615 2119
rect 67543 2079 67615 2085
rect 67543 2069 67575 2079
rect 67383 2017 67417 2069
rect 67549 2017 67575 2069
rect 67583 2069 67615 2079
rect 67743 2085 67775 2119
rect 67783 2085 67815 2119
rect 67743 2079 67815 2085
rect 67743 2069 67775 2079
rect 67583 2017 67617 2069
rect 67749 2017 67775 2069
rect 67783 2069 67815 2079
rect 67943 2085 67975 2119
rect 67983 2085 68015 2119
rect 67943 2079 68015 2085
rect 67943 2069 67975 2079
rect 67783 2017 67817 2069
rect 67949 2017 67975 2069
rect 67983 2069 68015 2079
rect 68143 2085 68175 2119
rect 68183 2085 68215 2119
rect 68143 2079 68215 2085
rect 68143 2069 68175 2079
rect 67983 2017 68017 2069
rect 68149 2017 68175 2069
rect 68183 2069 68215 2079
rect 68343 2069 68615 2119
rect 68743 2085 68775 2119
rect 68799 2085 68809 2119
rect 68743 2079 68811 2085
rect 68743 2069 68775 2079
rect 68183 2017 68217 2069
rect 68347 2017 68617 2069
rect 68764 2058 68775 2069
rect -53 1983 68879 2017
rect -53 1947 493 1983
rect 1147 1947 1411 1983
rect 3947 1947 4211 1983
rect 4747 1947 5011 1983
rect 8947 1947 9211 1983
rect 9347 1947 9611 1983
rect 10747 1947 11011 1983
rect 11147 1947 11411 1983
rect 12547 1947 12811 1983
rect 12947 1947 13211 1983
rect 14347 1947 14611 1983
rect 14747 1947 15011 1983
rect 16147 1947 16411 1983
rect 16547 1947 16811 1983
rect 19347 1947 19611 1983
rect 20147 1947 20411 1983
rect 21547 1947 21811 1983
rect 21947 1947 22211 1983
rect 23347 1947 23611 1983
rect 23747 1947 24011 1983
rect 25147 1947 25411 1983
rect 25547 1947 25811 1983
rect 26947 1947 27211 1983
rect 27347 1947 27611 1983
rect 28747 1947 29011 1983
rect 29147 1947 29411 1983
rect 30547 1947 30811 1983
rect 30947 1947 31211 1983
rect 32347 1947 32611 1983
rect 32747 1947 33011 1983
rect 34147 1947 34411 1983
rect 34547 1947 34811 1983
rect 35947 1947 36211 1983
rect 36347 1947 36611 1983
rect 37747 1947 38011 1983
rect 38147 1947 38411 1983
rect 39547 1947 39811 1983
rect 39947 1947 40211 1983
rect 41347 1947 41611 1983
rect 41747 1947 42011 1983
rect 43147 1947 43411 1983
rect 43547 1947 43811 1983
rect 44947 1947 45211 1983
rect 45347 1947 45611 1983
rect 46747 1947 47011 1983
rect 47147 1947 47411 1983
rect 48547 1947 48811 1983
rect 48947 1947 49211 1983
rect 50347 1947 50611 1983
rect 50747 1947 51011 1983
rect 52147 1947 52411 1983
rect 52547 1947 52811 1983
rect 53947 1947 54211 1983
rect 54347 1947 54611 1983
rect 55747 1947 56011 1983
rect 56147 1947 56411 1983
rect 57547 1947 57811 1983
rect 57947 1947 58211 1983
rect 59347 1947 59611 1983
rect 59747 1947 60011 1983
rect 61147 1947 61411 1983
rect 61547 1947 61811 1983
rect 62947 1947 63211 1983
rect 63347 1947 63611 1983
rect 64747 1947 65011 1983
rect 65147 1947 65411 1983
rect 66547 1947 66811 1983
rect 66947 1947 67211 1983
rect 68347 1947 68611 1983
rect -52 1747 489 1947
rect -52 1713 1355 1747
rect -52 1661 488 1713
rect 541 1679 547 1713
rect 741 1679 747 1713
rect 941 1679 947 1713
rect 1141 1679 1147 1713
rect 525 1661 583 1679
rect 725 1661 783 1679
rect 925 1661 983 1679
rect 1125 1661 1196 1679
rect 1199 1661 1251 1679
rect -52 1651 491 1661
rect 525 1651 691 1661
rect 725 1651 891 1661
rect 925 1651 1091 1661
rect -52 1561 493 1651
rect 525 1645 693 1651
rect 725 1645 893 1651
rect 925 1645 1093 1651
rect 1125 1645 1251 1661
rect 541 1561 693 1645
rect 741 1561 893 1645
rect 941 1561 1093 1645
rect 1141 1611 1275 1645
rect 1141 1572 1251 1611
rect 1141 1561 1291 1572
rect 1307 1561 1337 1577
rect -52 1401 1337 1561
rect 1341 1401 1451 1651
rect -53 1357 1451 1401
rect 4747 1365 4812 1383
rect 9347 1365 9412 1383
rect 11147 1365 11212 1383
rect 12947 1365 13012 1383
rect 14747 1365 14812 1383
rect 16547 1365 16612 1383
rect 20147 1365 20212 1383
rect 21947 1365 22012 1383
rect 23747 1365 23812 1383
rect 25547 1365 25612 1383
rect 27347 1365 27412 1383
rect 29147 1365 29212 1383
rect 30947 1365 31012 1383
rect 32747 1365 32812 1383
rect 34547 1365 34612 1383
rect 36347 1365 36412 1383
rect 38147 1365 38212 1383
rect 39947 1365 40012 1383
rect 41747 1365 41812 1383
rect 43547 1365 43612 1383
rect 45347 1365 45412 1383
rect 47147 1365 47212 1383
rect 48947 1365 49012 1383
rect 50747 1365 50812 1383
rect 52547 1365 52612 1383
rect 54347 1365 54412 1383
rect 56147 1365 56212 1383
rect 57947 1365 58012 1383
rect 59747 1365 59812 1383
rect 61547 1365 61612 1383
rect 63347 1365 63412 1383
rect 65147 1365 65212 1383
rect 66947 1365 67012 1383
rect -53 1353 1337 1357
rect -53 1347 1251 1353
rect 1341 1347 1451 1357
rect -53 1313 1485 1347
rect 2679 1313 2885 1347
rect 4079 1331 4280 1365
rect -53 1285 1275 1313
rect -53 1269 1251 1285
rect -53 1251 1212 1269
rect 1240 1258 1251 1269
rect -53 1217 1223 1251
rect 1341 1245 1451 1313
rect 4349 1269 4376 1365
rect 1343 1227 1451 1245
rect 1341 1217 1451 1227
rect -53 1183 1451 1217
rect -53 1147 1223 1183
rect 1297 1173 1337 1177
rect 1427 1173 1467 1177
rect 1285 1172 1343 1173
rect 1421 1172 1467 1173
rect 1285 1158 1348 1172
rect 1416 1161 1467 1172
rect 1421 1158 1467 1161
rect -17 879 18 1147
rect 97 978 132 1147
rect 227 978 262 1147
rect 159 885 200 919
rect 341 879 376 1147
rect 349 819 376 879
rect -17 817 18 819
rect 341 817 376 819
rect -17 783 376 817
rect 383 817 418 1147
rect 497 978 532 1147
rect 627 978 662 1147
rect 547 919 612 925
rect 547 885 600 919
rect 547 879 612 885
rect 741 879 776 1147
rect 749 819 776 879
rect 741 817 776 819
rect 383 783 776 817
rect 783 817 818 1147
rect 897 978 932 1147
rect 1027 978 1062 1147
rect 947 919 1012 925
rect 947 885 1000 919
rect 947 879 1012 885
rect 1141 879 1223 1147
rect 1297 969 1337 1158
rect 1343 969 1348 1158
rect 1427 969 1467 1158
rect 1347 919 1417 925
rect 1347 885 1405 919
rect 1347 879 1417 885
rect 1541 879 1581 1251
rect 2583 879 2623 1251
rect 2759 1211 2805 1245
rect 2697 969 2737 1161
rect 2743 969 2748 1172
rect 2816 1161 2821 1172
rect 2827 969 2867 1161
rect 2747 919 2817 925
rect 2747 885 2805 919
rect 2747 879 2817 885
rect 2941 879 2981 1251
rect 3983 879 4018 1269
rect 4159 1229 4200 1263
rect 4097 978 4132 1170
rect 4227 978 4262 1170
rect 4147 919 4212 925
rect 4147 885 4200 919
rect 4147 879 4212 885
rect 4341 879 4376 1269
rect 1147 819 1223 879
rect 4349 819 4376 879
rect 1141 817 1223 819
rect 3983 817 4018 819
rect 4341 817 4376 819
rect 783 801 1230 817
rect 1279 801 1485 817
rect 2679 801 2885 817
rect 783 783 1581 801
rect 2583 783 2981 801
rect 3983 783 4376 817
rect 4383 1331 4430 1365
rect 4479 1331 4680 1365
rect 4729 1347 4812 1365
rect 4383 817 4418 1331
rect 4747 1313 4830 1347
rect 4879 1313 5085 1347
rect 6279 1313 6485 1347
rect 7679 1313 7885 1347
rect 9079 1331 9280 1365
rect 9329 1347 9412 1365
rect 9347 1313 9430 1347
rect 9479 1313 9685 1347
rect 10879 1331 11080 1365
rect 11129 1347 11212 1365
rect 11147 1313 11230 1347
rect 11279 1313 11485 1347
rect 12679 1331 12880 1365
rect 12929 1347 13012 1365
rect 12947 1313 13030 1347
rect 13079 1313 13285 1347
rect 14479 1331 14680 1365
rect 14729 1347 14812 1365
rect 14747 1313 14830 1347
rect 14879 1313 15085 1347
rect 16279 1331 16480 1365
rect 16529 1347 16612 1365
rect 16547 1313 16630 1347
rect 16679 1313 16885 1347
rect 18079 1313 18285 1347
rect 19479 1331 19680 1365
rect 4747 1269 4823 1313
rect 9347 1269 9423 1313
rect 11147 1269 11223 1313
rect 12947 1269 13023 1313
rect 14747 1269 14823 1313
rect 16547 1269 16623 1313
rect 19749 1269 19776 1365
rect 4559 1229 4600 1263
rect 4497 978 4532 1170
rect 4627 978 4662 1170
rect 4547 919 4612 925
rect 4547 885 4600 919
rect 4547 879 4612 885
rect 4741 879 4823 1269
rect 4959 1211 5005 1245
rect 4897 969 4937 1161
rect 4943 969 4948 1172
rect 5016 1161 5021 1172
rect 5027 969 5067 1161
rect 4947 919 5017 925
rect 4947 885 5005 919
rect 4947 879 5017 885
rect 5141 879 5181 1251
rect 6183 879 6223 1251
rect 6359 1211 6405 1245
rect 6297 969 6337 1161
rect 6343 969 6348 1172
rect 6416 1161 6421 1172
rect 6427 969 6467 1161
rect 6347 919 6417 925
rect 6347 885 6405 919
rect 6347 879 6417 885
rect 6541 879 6581 1251
rect 7583 879 7623 1251
rect 7759 1211 7805 1245
rect 7697 969 7737 1161
rect 7743 969 7748 1172
rect 7816 1161 7821 1172
rect 7827 969 7867 1161
rect 7747 919 7817 925
rect 7747 885 7805 919
rect 7747 879 7817 885
rect 7941 879 7981 1251
rect 8983 879 9018 1269
rect 9159 1229 9200 1263
rect 9097 978 9132 1170
rect 9227 978 9262 1170
rect 9147 919 9212 925
rect 9147 885 9200 919
rect 9147 879 9212 885
rect 9341 879 9423 1269
rect 9559 1211 9605 1245
rect 9497 969 9537 1161
rect 9543 969 9548 1172
rect 9616 1161 9621 1172
rect 9627 969 9667 1161
rect 9547 919 9617 925
rect 9547 885 9605 919
rect 9547 879 9617 885
rect 9741 879 9781 1251
rect 10783 879 10818 1269
rect 10959 1229 11000 1263
rect 10897 978 10932 1170
rect 11027 978 11062 1170
rect 10947 919 11012 925
rect 10947 885 11000 919
rect 10947 879 11012 885
rect 11141 879 11223 1269
rect 11359 1211 11405 1245
rect 11297 969 11337 1161
rect 11343 969 11348 1172
rect 11416 1161 11421 1172
rect 11427 969 11467 1161
rect 11347 919 11417 925
rect 11347 885 11405 919
rect 11347 879 11417 885
rect 11541 879 11581 1251
rect 12583 879 12618 1269
rect 12759 1229 12800 1263
rect 12697 978 12732 1170
rect 12827 978 12862 1170
rect 12747 919 12812 925
rect 12747 885 12800 919
rect 12747 879 12812 885
rect 12941 879 13023 1269
rect 13159 1211 13205 1245
rect 13097 969 13137 1161
rect 13143 969 13148 1172
rect 13216 1161 13221 1172
rect 13227 969 13267 1161
rect 13147 919 13217 925
rect 13147 885 13205 919
rect 13147 879 13217 885
rect 13341 879 13381 1251
rect 14383 879 14418 1269
rect 14559 1229 14600 1263
rect 14497 978 14532 1170
rect 14627 978 14662 1170
rect 14547 919 14612 925
rect 14547 885 14600 919
rect 14547 879 14612 885
rect 14741 879 14823 1269
rect 14959 1211 15005 1245
rect 14897 969 14937 1161
rect 14943 969 14948 1172
rect 15016 1161 15021 1172
rect 15027 969 15067 1161
rect 14947 919 15017 925
rect 14947 885 15005 919
rect 14947 879 15017 885
rect 15141 879 15181 1251
rect 16183 879 16218 1269
rect 16347 1263 16412 1269
rect 16347 1229 16400 1263
rect 16347 1223 16412 1229
rect 16319 1195 16440 1200
rect 16297 978 16332 1170
rect 16427 978 16462 1170
rect 16347 919 16412 925
rect 16347 885 16400 919
rect 16347 879 16412 885
rect 16541 879 16623 1269
rect 16747 1245 16817 1251
rect 16747 1228 16805 1245
rect 16747 1205 16817 1228
rect 16719 1177 16845 1200
rect 16697 969 16737 1161
rect 16743 969 16748 1172
rect 16816 1161 16821 1172
rect 16827 969 16867 1161
rect 16747 919 16817 925
rect 16747 885 16805 919
rect 16747 879 16817 885
rect 16941 879 16981 1251
rect 17983 879 18023 1251
rect 18147 1245 18217 1251
rect 18147 1228 18205 1245
rect 18147 1205 18217 1228
rect 18119 1177 18245 1200
rect 18097 969 18137 1161
rect 18143 969 18148 1172
rect 18216 1161 18221 1172
rect 18227 969 18267 1161
rect 18147 919 18217 925
rect 18147 885 18205 919
rect 18147 879 18217 885
rect 18341 879 18381 1251
rect 19383 879 19418 1269
rect 19547 1263 19612 1269
rect 19547 1229 19600 1263
rect 19547 1223 19612 1229
rect 19519 1195 19640 1200
rect 19497 978 19532 1170
rect 19627 978 19662 1170
rect 19547 919 19612 925
rect 19547 885 19600 919
rect 19547 879 19612 885
rect 19741 879 19776 1269
rect 4747 819 4823 879
rect 9347 819 9423 879
rect 11147 819 11223 879
rect 12947 819 13023 879
rect 14747 819 14823 879
rect 16547 819 16623 879
rect 19749 819 19776 879
rect 4741 817 4823 819
rect 8983 817 9018 819
rect 9341 817 9423 819
rect 10783 817 10818 819
rect 11141 817 11223 819
rect 12583 817 12618 819
rect 12941 817 13023 819
rect 14383 817 14418 819
rect 14741 817 14823 819
rect 16183 817 16218 819
rect 16541 817 16623 819
rect 19383 817 19418 819
rect 19741 817 19776 819
rect 4383 801 4830 817
rect 4879 801 5085 817
rect 6279 801 6485 817
rect 7679 801 7885 817
rect 8983 801 9430 817
rect 9479 801 9685 817
rect 10783 801 11230 817
rect 11279 801 11485 817
rect 12583 801 13030 817
rect 13079 801 13285 817
rect 14383 801 14830 817
rect 14879 801 15085 817
rect 16183 801 16630 817
rect 16679 801 16885 817
rect 18079 801 18285 817
rect 4383 783 5181 801
rect 6183 783 6581 801
rect 7583 783 7981 801
rect 8983 783 9781 801
rect 10783 783 11581 801
rect 12583 783 13381 801
rect 14383 783 15181 801
rect 16183 783 16981 801
rect 17983 783 18381 801
rect 19383 783 19776 817
rect 19783 1331 19830 1365
rect 19879 1331 20080 1365
rect 20129 1347 20212 1365
rect 19783 817 19818 1331
rect 20147 1313 20230 1347
rect 20279 1313 20485 1347
rect 21679 1331 21880 1365
rect 21929 1347 22012 1365
rect 21947 1313 22030 1347
rect 22079 1313 22285 1347
rect 23479 1331 23680 1365
rect 23729 1347 23812 1365
rect 23747 1313 23830 1347
rect 23879 1313 24085 1347
rect 25279 1331 25480 1365
rect 25529 1347 25612 1365
rect 25547 1313 25630 1347
rect 25679 1313 25885 1347
rect 27079 1331 27280 1365
rect 27329 1347 27412 1365
rect 27347 1313 27430 1347
rect 27479 1313 27685 1347
rect 28879 1331 29080 1365
rect 29129 1347 29212 1365
rect 29147 1313 29230 1347
rect 29279 1313 29485 1347
rect 30679 1331 30880 1365
rect 30929 1347 31012 1365
rect 30947 1313 31030 1347
rect 31079 1313 31285 1347
rect 32479 1331 32680 1365
rect 32729 1347 32812 1365
rect 32747 1313 32830 1347
rect 32879 1313 33085 1347
rect 34279 1331 34480 1365
rect 34529 1347 34612 1365
rect 34547 1313 34630 1347
rect 34679 1313 34885 1347
rect 36079 1331 36280 1365
rect 36329 1347 36412 1365
rect 36347 1313 36430 1347
rect 36479 1313 36685 1347
rect 37879 1331 38080 1365
rect 38129 1347 38212 1365
rect 38147 1313 38230 1347
rect 38279 1313 38485 1347
rect 39679 1331 39880 1365
rect 39929 1347 40012 1365
rect 39947 1313 40030 1347
rect 40079 1313 40285 1347
rect 41479 1331 41680 1365
rect 41729 1347 41812 1365
rect 41747 1313 41830 1347
rect 41879 1313 42085 1347
rect 43279 1331 43480 1365
rect 43529 1347 43612 1365
rect 43547 1313 43630 1347
rect 43679 1313 43885 1347
rect 45079 1331 45280 1365
rect 45329 1347 45412 1365
rect 45347 1313 45430 1347
rect 45479 1313 45685 1347
rect 46879 1331 47080 1365
rect 47129 1347 47212 1365
rect 47147 1313 47230 1347
rect 47279 1313 47485 1347
rect 48679 1331 48880 1365
rect 48929 1347 49012 1365
rect 48947 1313 49030 1347
rect 49079 1313 49285 1347
rect 50479 1331 50680 1365
rect 50729 1347 50812 1365
rect 50747 1313 50830 1347
rect 50879 1313 51085 1347
rect 52279 1331 52480 1365
rect 52529 1347 52612 1365
rect 52547 1313 52630 1347
rect 52679 1313 52885 1347
rect 54079 1331 54280 1365
rect 54329 1347 54412 1365
rect 54347 1313 54430 1347
rect 54479 1313 54685 1347
rect 55879 1331 56080 1365
rect 56129 1347 56212 1365
rect 56147 1313 56230 1347
rect 56279 1313 56485 1347
rect 57679 1331 57880 1365
rect 57929 1347 58012 1365
rect 57947 1313 58030 1347
rect 58079 1313 58285 1347
rect 59479 1331 59680 1365
rect 59729 1347 59812 1365
rect 59747 1313 59830 1347
rect 59879 1313 60085 1347
rect 61279 1331 61480 1365
rect 61529 1347 61612 1365
rect 61547 1313 61630 1347
rect 61679 1313 61885 1347
rect 63079 1331 63280 1365
rect 63329 1347 63412 1365
rect 63347 1313 63430 1347
rect 63479 1313 63685 1347
rect 64879 1331 65080 1365
rect 65129 1347 65212 1365
rect 65147 1313 65230 1347
rect 65279 1313 65485 1347
rect 66679 1331 66880 1365
rect 66929 1347 67012 1365
rect 66947 1313 67030 1347
rect 67079 1313 67285 1347
rect 68479 1331 68680 1365
rect 20147 1269 20223 1313
rect 21947 1269 22023 1313
rect 23747 1269 23823 1313
rect 25547 1269 25623 1313
rect 27347 1269 27423 1313
rect 29147 1269 29223 1313
rect 30947 1269 31023 1313
rect 32747 1269 32823 1313
rect 34547 1269 34623 1313
rect 36347 1269 36423 1313
rect 38147 1269 38223 1313
rect 39947 1269 40023 1313
rect 41747 1269 41823 1313
rect 43547 1269 43623 1313
rect 45347 1269 45423 1313
rect 47147 1269 47223 1313
rect 48947 1269 49023 1313
rect 50747 1269 50823 1313
rect 52547 1269 52623 1313
rect 54347 1269 54423 1313
rect 56147 1269 56223 1313
rect 57947 1269 58023 1313
rect 59747 1269 59823 1313
rect 61547 1269 61623 1313
rect 63347 1269 63423 1313
rect 65147 1269 65223 1313
rect 66947 1269 67023 1313
rect 19947 1263 20012 1269
rect 19947 1229 20000 1263
rect 19947 1223 20012 1229
rect 19919 1195 20040 1200
rect 19897 978 19932 1170
rect 20027 978 20062 1170
rect 19947 919 20012 925
rect 19947 885 20000 919
rect 19947 879 20012 885
rect 20141 879 20223 1269
rect 20347 1245 20417 1251
rect 20347 1228 20405 1245
rect 20347 1205 20417 1228
rect 20319 1177 20445 1200
rect 20297 969 20337 1161
rect 20343 969 20348 1172
rect 20416 1161 20421 1172
rect 20427 969 20467 1161
rect 20347 919 20417 925
rect 20347 885 20405 919
rect 20347 879 20417 885
rect 20541 879 20581 1251
rect 21583 879 21618 1269
rect 21747 1263 21812 1269
rect 21747 1229 21800 1263
rect 21747 1223 21812 1229
rect 21719 1195 21840 1200
rect 21697 978 21732 1170
rect 21827 978 21862 1170
rect 21747 919 21812 925
rect 21747 885 21800 919
rect 21747 879 21812 885
rect 21941 879 22023 1269
rect 22147 1245 22217 1251
rect 22147 1228 22205 1245
rect 22147 1205 22217 1228
rect 22119 1177 22245 1200
rect 22097 969 22137 1161
rect 22143 969 22148 1172
rect 22216 1161 22221 1172
rect 22227 969 22267 1161
rect 22147 919 22217 925
rect 22147 885 22205 919
rect 22147 879 22217 885
rect 22341 879 22381 1251
rect 23383 879 23418 1269
rect 23547 1263 23612 1269
rect 23547 1229 23600 1263
rect 23547 1223 23612 1229
rect 23519 1195 23640 1200
rect 23497 978 23532 1170
rect 23627 978 23662 1170
rect 23547 919 23612 925
rect 23547 885 23600 919
rect 23547 879 23612 885
rect 23741 879 23823 1269
rect 23947 1245 24017 1251
rect 23947 1228 24005 1245
rect 23947 1205 24017 1228
rect 23919 1177 24045 1200
rect 23897 969 23937 1161
rect 23943 969 23948 1172
rect 24016 1161 24021 1172
rect 24027 969 24067 1161
rect 23947 919 24017 925
rect 23947 885 24005 919
rect 23947 879 24017 885
rect 24141 879 24181 1251
rect 25183 879 25218 1269
rect 25347 1263 25412 1269
rect 25347 1229 25400 1263
rect 25347 1223 25412 1229
rect 25319 1195 25440 1200
rect 25297 978 25332 1170
rect 25427 978 25462 1170
rect 25347 919 25412 925
rect 25347 885 25400 919
rect 25347 879 25412 885
rect 25541 879 25623 1269
rect 25747 1245 25817 1251
rect 25747 1228 25805 1245
rect 25747 1205 25817 1228
rect 25719 1177 25845 1200
rect 25697 969 25737 1161
rect 25743 969 25748 1172
rect 25816 1161 25821 1172
rect 25827 969 25867 1161
rect 25747 919 25817 925
rect 25747 885 25805 919
rect 25747 879 25817 885
rect 25941 879 25981 1251
rect 26983 879 27018 1269
rect 27147 1263 27212 1269
rect 27147 1229 27200 1263
rect 27147 1223 27212 1229
rect 27119 1195 27240 1200
rect 27097 978 27132 1170
rect 27227 978 27262 1170
rect 27147 919 27212 925
rect 27147 885 27200 919
rect 27147 879 27212 885
rect 27341 879 27423 1269
rect 27547 1245 27617 1251
rect 27547 1228 27605 1245
rect 27547 1205 27617 1228
rect 27519 1177 27645 1200
rect 27497 969 27537 1161
rect 27543 969 27548 1172
rect 27616 1161 27621 1172
rect 27627 969 27667 1161
rect 27547 919 27617 925
rect 27547 885 27605 919
rect 27547 879 27617 885
rect 27741 879 27781 1251
rect 28783 879 28818 1269
rect 28947 1263 29012 1269
rect 28947 1229 29000 1263
rect 28947 1223 29012 1229
rect 28919 1195 29040 1200
rect 28897 978 28932 1170
rect 29027 978 29062 1170
rect 28947 919 29012 925
rect 28947 885 29000 919
rect 28947 879 29012 885
rect 29141 879 29223 1269
rect 29347 1245 29417 1251
rect 29347 1228 29405 1245
rect 29347 1205 29417 1228
rect 29319 1177 29445 1200
rect 29297 969 29337 1161
rect 29343 969 29348 1172
rect 29416 1161 29421 1172
rect 29427 969 29467 1161
rect 29347 919 29417 925
rect 29347 885 29405 919
rect 29347 879 29417 885
rect 29541 879 29581 1251
rect 30583 879 30618 1269
rect 30747 1263 30812 1269
rect 30747 1229 30800 1263
rect 30747 1223 30812 1229
rect 30719 1195 30840 1200
rect 30697 978 30732 1170
rect 30827 978 30862 1170
rect 30747 919 30812 925
rect 30747 885 30800 919
rect 30747 879 30812 885
rect 30941 879 31023 1269
rect 31147 1245 31217 1251
rect 31147 1228 31205 1245
rect 31147 1205 31217 1228
rect 31119 1177 31245 1200
rect 31097 969 31137 1161
rect 31143 969 31148 1172
rect 31216 1161 31221 1172
rect 31227 969 31267 1161
rect 31147 919 31217 925
rect 31147 885 31205 919
rect 31147 879 31217 885
rect 31341 879 31381 1251
rect 32383 879 32418 1269
rect 32547 1263 32612 1269
rect 32547 1229 32600 1263
rect 32547 1223 32612 1229
rect 32519 1195 32640 1200
rect 32497 978 32532 1170
rect 32627 978 32662 1170
rect 32547 919 32612 925
rect 32547 885 32600 919
rect 32547 879 32612 885
rect 32741 879 32823 1269
rect 32947 1245 33017 1251
rect 32947 1228 33005 1245
rect 32947 1205 33017 1228
rect 32919 1177 33045 1200
rect 32897 969 32937 1161
rect 32943 969 32948 1172
rect 33016 1161 33021 1172
rect 33027 969 33067 1161
rect 32947 919 33017 925
rect 32947 885 33005 919
rect 32947 879 33017 885
rect 33141 879 33181 1251
rect 34183 879 34218 1269
rect 34347 1263 34412 1269
rect 34347 1229 34400 1263
rect 34347 1223 34412 1229
rect 34319 1195 34440 1200
rect 34297 978 34332 1170
rect 34427 978 34462 1170
rect 34347 919 34412 925
rect 34347 885 34400 919
rect 34347 879 34412 885
rect 34541 879 34623 1269
rect 34747 1245 34817 1251
rect 34747 1228 34805 1245
rect 34747 1205 34817 1228
rect 34719 1177 34845 1200
rect 34697 969 34737 1161
rect 34743 969 34748 1172
rect 34816 1161 34821 1172
rect 34827 969 34867 1161
rect 34747 919 34817 925
rect 34747 885 34805 919
rect 34747 879 34817 885
rect 34941 879 34981 1251
rect 35983 879 36018 1269
rect 36147 1263 36212 1269
rect 36147 1229 36200 1263
rect 36147 1223 36212 1229
rect 36119 1195 36240 1200
rect 36097 978 36132 1170
rect 36227 978 36262 1170
rect 36147 919 36212 925
rect 36147 885 36200 919
rect 36147 879 36212 885
rect 36341 879 36423 1269
rect 36547 1245 36617 1251
rect 36547 1228 36605 1245
rect 36547 1205 36617 1228
rect 36519 1177 36645 1200
rect 36497 969 36537 1161
rect 36543 969 36548 1172
rect 36616 1161 36621 1172
rect 36627 969 36667 1161
rect 36547 919 36617 925
rect 36547 885 36605 919
rect 36547 879 36617 885
rect 36741 879 36781 1251
rect 37783 879 37818 1269
rect 37947 1263 38012 1269
rect 37947 1229 38000 1263
rect 37947 1223 38012 1229
rect 37919 1195 38040 1200
rect 37897 978 37932 1170
rect 38027 978 38062 1170
rect 37947 919 38012 925
rect 37947 885 38000 919
rect 37947 879 38012 885
rect 38141 879 38223 1269
rect 38347 1245 38417 1251
rect 38347 1228 38405 1245
rect 38347 1205 38417 1228
rect 38319 1177 38445 1200
rect 38297 969 38337 1161
rect 38343 969 38348 1172
rect 38416 1161 38421 1172
rect 38427 969 38467 1161
rect 38347 919 38417 925
rect 38347 885 38405 919
rect 38347 879 38417 885
rect 38541 879 38581 1251
rect 39583 879 39618 1269
rect 39747 1263 39812 1269
rect 39747 1229 39800 1263
rect 39747 1223 39812 1229
rect 39719 1195 39840 1200
rect 39697 978 39732 1170
rect 39827 978 39862 1170
rect 39747 919 39812 925
rect 39747 885 39800 919
rect 39747 879 39812 885
rect 39941 879 40023 1269
rect 40147 1245 40217 1251
rect 40147 1228 40205 1245
rect 40147 1205 40217 1228
rect 40119 1177 40245 1200
rect 40097 969 40137 1161
rect 40143 969 40148 1172
rect 40216 1161 40221 1172
rect 40227 969 40267 1161
rect 40147 919 40217 925
rect 40147 885 40205 919
rect 40147 879 40217 885
rect 40341 879 40381 1251
rect 41383 879 41418 1269
rect 41547 1263 41612 1269
rect 41547 1229 41600 1263
rect 41547 1223 41612 1229
rect 41519 1195 41640 1200
rect 41497 978 41532 1170
rect 41627 978 41662 1170
rect 41547 919 41612 925
rect 41547 885 41600 919
rect 41547 879 41612 885
rect 41741 879 41823 1269
rect 41947 1245 42017 1251
rect 41947 1228 42005 1245
rect 41947 1205 42017 1228
rect 41919 1177 42045 1200
rect 41897 969 41937 1161
rect 41943 969 41948 1172
rect 42016 1161 42021 1172
rect 42027 969 42067 1161
rect 41947 919 42017 925
rect 41947 885 42005 919
rect 41947 879 42017 885
rect 42141 879 42181 1251
rect 43183 879 43218 1269
rect 43347 1263 43412 1269
rect 43347 1229 43400 1263
rect 43347 1223 43412 1229
rect 43319 1195 43440 1200
rect 43297 978 43332 1170
rect 43427 978 43462 1170
rect 43347 919 43412 925
rect 43347 885 43400 919
rect 43347 879 43412 885
rect 43541 879 43623 1269
rect 43747 1245 43817 1251
rect 43747 1228 43805 1245
rect 43747 1205 43817 1228
rect 43719 1177 43845 1200
rect 43697 969 43737 1161
rect 43743 969 43748 1172
rect 43816 1161 43821 1172
rect 43827 969 43867 1161
rect 43747 919 43817 925
rect 43747 885 43805 919
rect 43747 879 43817 885
rect 43941 879 43981 1251
rect 44983 879 45018 1269
rect 45147 1263 45212 1269
rect 45147 1229 45200 1263
rect 45147 1223 45212 1229
rect 45119 1195 45240 1200
rect 45097 978 45132 1170
rect 45227 978 45262 1170
rect 45147 919 45212 925
rect 45147 885 45200 919
rect 45147 879 45212 885
rect 45341 879 45423 1269
rect 45547 1245 45617 1251
rect 45547 1228 45605 1245
rect 45547 1205 45617 1228
rect 45519 1177 45645 1200
rect 45497 969 45537 1161
rect 45543 969 45548 1172
rect 45616 1161 45621 1172
rect 45627 969 45667 1161
rect 45547 919 45617 925
rect 45547 885 45605 919
rect 45547 879 45617 885
rect 45741 879 45781 1251
rect 46783 879 46818 1269
rect 46947 1263 47012 1269
rect 46947 1229 47000 1263
rect 46947 1223 47012 1229
rect 46919 1195 47040 1200
rect 46897 978 46932 1170
rect 47027 978 47062 1170
rect 46947 919 47012 925
rect 46947 885 47000 919
rect 46947 879 47012 885
rect 47141 879 47223 1269
rect 47347 1245 47417 1251
rect 47347 1228 47405 1245
rect 47347 1205 47417 1228
rect 47319 1177 47445 1200
rect 47297 969 47337 1161
rect 47343 969 47348 1172
rect 47416 1161 47421 1172
rect 47427 969 47467 1161
rect 47347 919 47417 925
rect 47347 885 47405 919
rect 47347 879 47417 885
rect 47541 879 47581 1251
rect 48583 879 48618 1269
rect 48747 1263 48812 1269
rect 48747 1229 48800 1263
rect 48747 1223 48812 1229
rect 48719 1195 48840 1200
rect 48697 978 48732 1170
rect 48827 978 48862 1170
rect 48747 919 48812 925
rect 48747 885 48800 919
rect 48747 879 48812 885
rect 48941 879 49023 1269
rect 49147 1245 49217 1251
rect 49147 1228 49205 1245
rect 49147 1205 49217 1228
rect 49119 1177 49245 1200
rect 49097 969 49137 1161
rect 49143 969 49148 1172
rect 49216 1161 49221 1172
rect 49227 969 49267 1161
rect 49147 919 49217 925
rect 49147 885 49205 919
rect 49147 879 49217 885
rect 49341 879 49381 1251
rect 50383 879 50418 1269
rect 50547 1263 50612 1269
rect 50547 1229 50600 1263
rect 50547 1223 50612 1229
rect 50519 1195 50640 1200
rect 50497 978 50532 1170
rect 50627 978 50662 1170
rect 50547 919 50612 925
rect 50547 885 50600 919
rect 50547 879 50612 885
rect 50741 879 50823 1269
rect 50947 1245 51017 1251
rect 50947 1228 51005 1245
rect 50947 1205 51017 1228
rect 50919 1177 51045 1200
rect 50897 969 50937 1161
rect 50943 969 50948 1172
rect 51016 1161 51021 1172
rect 51027 969 51067 1161
rect 50947 919 51017 925
rect 50947 885 51005 919
rect 50947 879 51017 885
rect 51141 879 51181 1251
rect 52183 879 52218 1269
rect 52347 1263 52412 1269
rect 52347 1229 52400 1263
rect 52347 1223 52412 1229
rect 52319 1195 52440 1200
rect 52297 978 52332 1170
rect 52427 978 52462 1170
rect 52347 919 52412 925
rect 52347 885 52400 919
rect 52347 879 52412 885
rect 52541 879 52623 1269
rect 52747 1245 52817 1251
rect 52747 1228 52805 1245
rect 52747 1205 52817 1228
rect 52719 1177 52845 1200
rect 52697 969 52737 1161
rect 52743 969 52748 1172
rect 52816 1161 52821 1172
rect 52827 969 52867 1161
rect 52747 919 52817 925
rect 52747 885 52805 919
rect 52747 879 52817 885
rect 52941 879 52981 1251
rect 53983 879 54018 1269
rect 54147 1263 54212 1269
rect 54147 1229 54200 1263
rect 54147 1223 54212 1229
rect 54119 1195 54240 1200
rect 54097 978 54132 1170
rect 54227 978 54262 1170
rect 54147 919 54212 925
rect 54147 885 54200 919
rect 54147 879 54212 885
rect 54341 879 54423 1269
rect 54547 1245 54617 1251
rect 54547 1228 54605 1245
rect 54547 1205 54617 1228
rect 54519 1177 54645 1200
rect 54497 969 54537 1161
rect 54543 969 54548 1172
rect 54616 1161 54621 1172
rect 54627 969 54667 1161
rect 54547 919 54617 925
rect 54547 885 54605 919
rect 54547 879 54617 885
rect 54741 879 54781 1251
rect 55783 879 55818 1269
rect 55947 1263 56012 1269
rect 55947 1229 56000 1263
rect 55947 1223 56012 1229
rect 55919 1195 56040 1200
rect 55897 978 55932 1170
rect 56027 978 56062 1170
rect 55947 919 56012 925
rect 55947 885 56000 919
rect 55947 879 56012 885
rect 56141 879 56223 1269
rect 56347 1245 56417 1251
rect 56347 1228 56405 1245
rect 56347 1205 56417 1228
rect 56319 1177 56445 1200
rect 56297 969 56337 1161
rect 56343 969 56348 1172
rect 56416 1161 56421 1172
rect 56427 969 56467 1161
rect 56347 919 56417 925
rect 56347 885 56405 919
rect 56347 879 56417 885
rect 56541 879 56581 1251
rect 57583 879 57618 1269
rect 57747 1263 57812 1269
rect 57747 1229 57800 1263
rect 57747 1223 57812 1229
rect 57719 1195 57840 1200
rect 57697 978 57732 1170
rect 57827 978 57862 1170
rect 57747 919 57812 925
rect 57747 885 57800 919
rect 57747 879 57812 885
rect 57941 879 58023 1269
rect 58147 1245 58217 1251
rect 58147 1228 58205 1245
rect 58147 1205 58217 1228
rect 58119 1177 58245 1200
rect 58097 969 58137 1161
rect 58143 969 58148 1172
rect 58216 1161 58221 1172
rect 58227 969 58267 1161
rect 58147 919 58217 925
rect 58147 885 58205 919
rect 58147 879 58217 885
rect 58341 879 58381 1251
rect 59383 879 59418 1269
rect 59547 1263 59612 1269
rect 59547 1229 59600 1263
rect 59547 1223 59612 1229
rect 59519 1195 59640 1200
rect 59497 978 59532 1170
rect 59627 978 59662 1170
rect 59547 919 59612 925
rect 59547 885 59600 919
rect 59547 879 59612 885
rect 59741 879 59823 1269
rect 59947 1245 60017 1251
rect 59947 1228 60005 1245
rect 59947 1205 60017 1228
rect 59919 1177 60045 1200
rect 59897 969 59937 1161
rect 59943 969 59948 1172
rect 60016 1161 60021 1172
rect 60027 969 60067 1161
rect 59947 919 60017 925
rect 59947 885 60005 919
rect 59947 879 60017 885
rect 60141 879 60181 1251
rect 61183 879 61218 1269
rect 61347 1263 61412 1269
rect 61347 1229 61400 1263
rect 61347 1223 61412 1229
rect 61319 1195 61440 1200
rect 61297 978 61332 1170
rect 61427 978 61462 1170
rect 61347 919 61412 925
rect 61347 885 61400 919
rect 61347 879 61412 885
rect 61541 879 61623 1269
rect 61747 1245 61817 1251
rect 61747 1228 61805 1245
rect 61747 1205 61817 1228
rect 61719 1177 61845 1200
rect 61697 969 61737 1161
rect 61743 969 61748 1172
rect 61816 1161 61821 1172
rect 61827 969 61867 1161
rect 61747 919 61817 925
rect 61747 885 61805 919
rect 61747 879 61817 885
rect 61941 879 61981 1251
rect 62983 879 63018 1269
rect 63147 1263 63212 1269
rect 63147 1229 63200 1263
rect 63147 1223 63212 1229
rect 63119 1195 63240 1200
rect 63097 978 63132 1170
rect 63227 978 63262 1170
rect 63147 919 63212 925
rect 63147 885 63200 919
rect 63147 879 63212 885
rect 63341 879 63423 1269
rect 63547 1245 63617 1251
rect 63547 1228 63605 1245
rect 63547 1205 63617 1228
rect 63519 1177 63645 1200
rect 63497 969 63537 1161
rect 63543 969 63548 1172
rect 63616 1161 63621 1172
rect 63627 969 63667 1161
rect 63547 919 63617 925
rect 63547 885 63605 919
rect 63547 879 63617 885
rect 63741 879 63781 1251
rect 64783 879 64818 1269
rect 64947 1263 65012 1269
rect 64947 1229 65000 1263
rect 64947 1223 65012 1229
rect 64919 1195 65040 1200
rect 64897 978 64932 1170
rect 65027 978 65062 1170
rect 64947 919 65012 925
rect 64947 885 65000 919
rect 64947 879 65012 885
rect 65141 879 65223 1269
rect 65347 1245 65417 1251
rect 65347 1228 65405 1245
rect 65347 1205 65417 1228
rect 65319 1177 65445 1200
rect 65297 969 65337 1161
rect 65343 969 65348 1172
rect 65416 1161 65421 1172
rect 65427 969 65467 1161
rect 65347 919 65417 925
rect 65347 885 65405 919
rect 65347 879 65417 885
rect 65541 879 65581 1251
rect 66583 879 66618 1269
rect 66747 1263 66812 1269
rect 66747 1229 66800 1263
rect 66747 1223 66812 1229
rect 66719 1195 66840 1200
rect 66697 978 66732 1170
rect 66827 978 66862 1170
rect 66747 919 66812 925
rect 66747 885 66800 919
rect 66747 879 66812 885
rect 66941 879 67023 1269
rect 67147 1245 67217 1251
rect 67147 1228 67205 1245
rect 67147 1205 67217 1228
rect 67119 1177 67245 1200
rect 67097 969 67137 1161
rect 67143 969 67148 1172
rect 67216 1161 67221 1172
rect 67227 969 67267 1161
rect 67147 919 67217 925
rect 67147 885 67205 919
rect 67147 879 67217 885
rect 67341 879 67381 1251
rect 68383 879 68418 1269
rect 68547 1263 68612 1269
rect 68547 1229 68600 1263
rect 68547 1223 68612 1229
rect 68519 1195 68640 1200
rect 68497 978 68532 1170
rect 68627 978 68662 1170
rect 68547 919 68612 925
rect 68547 885 68600 919
rect 68547 879 68612 885
rect 68741 879 68776 1269
rect 20147 819 20223 879
rect 21947 819 22023 879
rect 23747 819 23823 879
rect 25547 819 25623 879
rect 27347 819 27423 879
rect 29147 819 29223 879
rect 30947 819 31023 879
rect 32747 819 32823 879
rect 34547 819 34623 879
rect 36347 819 36423 879
rect 38147 819 38223 879
rect 39947 819 40023 879
rect 41747 819 41823 879
rect 43547 819 43623 879
rect 45347 819 45423 879
rect 47147 819 47223 879
rect 48947 819 49023 879
rect 50747 819 50823 879
rect 52547 819 52623 879
rect 54347 819 54423 879
rect 56147 819 56223 879
rect 57947 819 58023 879
rect 59747 819 59823 879
rect 61547 819 61623 879
rect 63347 819 63423 879
rect 65147 819 65223 879
rect 66947 819 67023 879
rect 20141 817 20223 819
rect 21583 817 21618 819
rect 21941 817 22023 819
rect 23383 817 23418 819
rect 23741 817 23823 819
rect 25183 817 25218 819
rect 25541 817 25623 819
rect 26983 817 27018 819
rect 27341 817 27423 819
rect 28783 817 28818 819
rect 29141 817 29223 819
rect 30583 817 30618 819
rect 30941 817 31023 819
rect 32383 817 32418 819
rect 32741 817 32823 819
rect 34183 817 34218 819
rect 34541 817 34623 819
rect 35983 817 36018 819
rect 36341 817 36423 819
rect 37783 817 37818 819
rect 38141 817 38223 819
rect 39583 817 39618 819
rect 39941 817 40023 819
rect 41383 817 41418 819
rect 41741 817 41823 819
rect 43183 817 43218 819
rect 43541 817 43623 819
rect 44983 817 45018 819
rect 45341 817 45423 819
rect 46783 817 46818 819
rect 47141 817 47223 819
rect 48583 817 48618 819
rect 48941 817 49023 819
rect 50383 817 50418 819
rect 50741 817 50823 819
rect 52183 817 52218 819
rect 52541 817 52623 819
rect 53983 817 54018 819
rect 54341 817 54423 819
rect 55783 817 55818 819
rect 56141 817 56223 819
rect 57583 817 57618 819
rect 57941 817 58023 819
rect 59383 817 59418 819
rect 59741 817 59823 819
rect 61183 817 61218 819
rect 61541 817 61623 819
rect 62983 817 63018 819
rect 63341 817 63423 819
rect 64783 817 64818 819
rect 65141 817 65223 819
rect 66583 817 66618 819
rect 66941 817 67023 819
rect 68383 817 68418 819
rect 68741 817 68776 819
rect 19783 801 20230 817
rect 20279 801 20485 817
rect 21583 801 22030 817
rect 22079 801 22285 817
rect 23383 801 23830 817
rect 23879 801 24085 817
rect 25183 801 25630 817
rect 25679 801 25885 817
rect 26983 801 27430 817
rect 27479 801 27685 817
rect 28783 801 29230 817
rect 29279 801 29485 817
rect 30583 801 31030 817
rect 31079 801 31285 817
rect 32383 801 32830 817
rect 32879 801 33085 817
rect 34183 801 34630 817
rect 34679 801 34885 817
rect 35983 801 36430 817
rect 36479 801 36685 817
rect 37783 801 38230 817
rect 38279 801 38485 817
rect 39583 801 40030 817
rect 40079 801 40285 817
rect 41383 801 41830 817
rect 41879 801 42085 817
rect 43183 801 43630 817
rect 43679 801 43885 817
rect 44983 801 45430 817
rect 45479 801 45685 817
rect 46783 801 47230 817
rect 47279 801 47485 817
rect 48583 801 49030 817
rect 49079 801 49285 817
rect 50383 801 50830 817
rect 50879 801 51085 817
rect 52183 801 52630 817
rect 52679 801 52885 817
rect 53983 801 54430 817
rect 54479 801 54685 817
rect 55783 801 56230 817
rect 56279 801 56485 817
rect 57583 801 58030 817
rect 58079 801 58285 817
rect 59383 801 59830 817
rect 59879 801 60085 817
rect 61183 801 61630 817
rect 61679 801 61885 817
rect 62983 801 63430 817
rect 63479 801 63685 817
rect 64783 801 65230 817
rect 65279 801 65485 817
rect 66583 801 67030 817
rect 67079 801 67285 817
rect 19783 783 20581 801
rect 21583 783 22381 801
rect 23383 783 24181 801
rect 25183 783 25981 801
rect 26983 783 27781 801
rect 28783 783 29581 801
rect 30583 783 31381 801
rect 32383 783 33181 801
rect 34183 783 34981 801
rect 35983 783 36781 801
rect 37783 783 38581 801
rect 39583 783 40381 801
rect 41383 783 42181 801
rect 43183 783 43981 801
rect 44983 783 45781 801
rect 46783 783 47581 801
rect 48583 783 49381 801
rect 50383 783 51181 801
rect 52183 783 52981 801
rect 53983 783 54781 801
rect 55783 783 56581 801
rect 57583 783 58381 801
rect 59383 783 60181 801
rect 61183 783 61981 801
rect 62983 783 63781 801
rect 64783 783 65581 801
rect 66583 783 67381 801
rect 68383 783 68776 817
rect 1147 765 1212 783
rect -17 749 375 765
rect 349 183 375 749
rect 383 749 775 765
rect 383 731 429 749
rect 383 217 417 731
rect 463 600 565 610
rect 593 600 695 610
rect 491 572 537 582
rect 621 572 667 582
rect 383 183 429 217
rect 749 183 775 749
rect 783 749 1212 765
rect 783 731 829 749
rect 1129 747 1212 749
rect 3947 765 4011 783
rect 4747 765 4812 783
rect 3947 749 4375 765
rect 783 217 817 731
rect 1147 713 1229 747
rect 1279 713 2479 747
rect 863 600 965 610
rect 993 600 1095 610
rect 891 572 937 582
rect 1021 572 1067 582
rect 1147 217 1217 713
rect 1549 679 1575 713
rect 1383 661 1394 672
rect 1343 611 1359 645
rect 1383 611 1415 661
rect 1525 651 1575 679
rect 1525 645 1541 651
rect 1543 611 1575 651
rect 1383 601 1417 611
rect 1541 601 1575 611
rect 1263 600 1365 601
rect 1383 600 1575 601
rect 1291 572 1337 573
rect 1383 319 1417 600
rect 1427 573 1451 577
rect 1507 573 1531 577
rect 1421 572 1467 573
rect 1427 353 1451 572
rect 1459 369 1461 561
rect 1463 400 1467 572
rect 1485 572 1537 573
rect 1485 357 1531 572
rect 1507 353 1531 357
rect 1541 353 1575 600
rect 1525 319 1575 353
rect 1343 285 1359 319
rect 1383 269 1415 319
rect 1543 269 1575 319
rect 1383 258 1394 269
rect 1549 217 1575 269
rect 1583 661 1617 713
rect 1749 679 1775 713
rect 1583 611 1615 661
rect 1725 651 1775 679
rect 1725 645 1741 651
rect 1743 611 1775 651
rect 1583 601 1617 611
rect 1741 601 1775 611
rect 1583 600 1775 601
rect 1583 319 1617 600
rect 1627 573 1651 577
rect 1707 573 1731 577
rect 1621 572 1667 573
rect 1627 353 1651 572
rect 1659 369 1661 561
rect 1663 400 1667 572
rect 1685 572 1737 573
rect 1685 357 1731 572
rect 1707 353 1731 357
rect 1741 353 1775 600
rect 1725 319 1775 353
rect 1583 269 1615 319
rect 1743 269 1775 319
rect 1583 217 1617 269
rect 1749 217 1775 269
rect 1783 661 1817 713
rect 1949 679 1975 713
rect 1783 611 1815 661
rect 1925 651 1975 679
rect 1925 645 1941 651
rect 1943 611 1975 651
rect 1783 601 1817 611
rect 1941 601 1975 611
rect 1783 600 1975 601
rect 1783 319 1817 600
rect 1827 573 1851 577
rect 1907 573 1931 577
rect 1821 572 1867 573
rect 1827 353 1851 572
rect 1859 369 1861 561
rect 1863 400 1867 572
rect 1885 572 1937 573
rect 1885 357 1931 572
rect 1907 353 1931 357
rect 1941 353 1975 600
rect 1925 319 1975 353
rect 1783 269 1815 319
rect 1943 269 1975 319
rect 1783 217 1817 269
rect 1949 217 1975 269
rect 1983 661 2017 713
rect 2149 679 2175 713
rect 1983 611 2015 661
rect 2125 651 2175 679
rect 2125 645 2141 651
rect 2143 611 2175 651
rect 1983 601 2017 611
rect 2141 601 2175 611
rect 1983 600 2175 601
rect 1983 319 2017 600
rect 2027 573 2051 577
rect 2107 573 2131 577
rect 2021 572 2067 573
rect 2027 353 2051 572
rect 2059 369 2061 561
rect 2063 400 2067 572
rect 2085 572 2137 573
rect 2085 357 2131 572
rect 2107 353 2131 357
rect 2141 353 2175 600
rect 2125 319 2175 353
rect 1983 269 2015 319
rect 2143 269 2175 319
rect 1983 217 2017 269
rect 2149 217 2175 269
rect 2183 661 2217 713
rect 2183 611 2215 661
rect 2325 651 2375 679
rect 2325 645 2341 651
rect 2343 611 2375 651
rect 2399 611 2409 645
rect 2183 601 2217 611
rect 2341 601 2375 611
rect 2183 600 2375 601
rect 2393 600 2495 601
rect 2183 319 2217 600
rect 2227 573 2251 577
rect 2307 573 2331 577
rect 2221 572 2267 573
rect 2227 353 2251 572
rect 2259 369 2261 561
rect 2263 400 2267 572
rect 2285 572 2337 573
rect 2285 357 2331 572
rect 2307 353 2331 357
rect 2341 353 2375 600
rect 2421 572 2467 573
rect 2325 319 2375 353
rect 2183 269 2215 319
rect 2343 269 2375 319
rect 2399 285 2409 319
rect 2183 217 2217 269
rect 2364 258 2375 269
rect 783 183 829 217
rect 1147 183 1229 217
rect 1279 183 2479 217
rect 2549 183 2575 747
rect 2583 713 2629 747
rect 2679 713 3879 747
rect 3947 731 4029 749
rect 2583 217 2617 713
rect 2949 679 2975 713
rect 2783 661 2794 672
rect 2743 611 2759 645
rect 2783 611 2815 661
rect 2925 651 2975 679
rect 2925 645 2941 651
rect 2943 611 2975 651
rect 2783 601 2817 611
rect 2941 601 2975 611
rect 2663 600 2765 601
rect 2783 600 2975 601
rect 2691 572 2737 573
rect 2783 319 2817 600
rect 2827 573 2851 577
rect 2907 573 2931 577
rect 2821 572 2867 573
rect 2827 353 2851 572
rect 2859 369 2861 561
rect 2863 400 2867 572
rect 2885 572 2937 573
rect 2885 357 2931 572
rect 2907 353 2931 357
rect 2941 353 2975 600
rect 2925 319 2975 353
rect 2743 285 2759 319
rect 2783 269 2815 319
rect 2943 269 2975 319
rect 2783 258 2794 269
rect 2949 217 2975 269
rect 2983 661 3017 713
rect 3149 679 3175 713
rect 2983 611 3015 661
rect 3125 651 3175 679
rect 3125 645 3141 651
rect 3143 611 3175 651
rect 2983 601 3017 611
rect 3141 601 3175 611
rect 2983 600 3175 601
rect 2983 319 3017 600
rect 3027 573 3051 577
rect 3107 573 3131 577
rect 3021 572 3067 573
rect 3027 353 3051 572
rect 3059 369 3061 561
rect 3063 400 3067 572
rect 3085 572 3137 573
rect 3085 357 3131 572
rect 3107 353 3131 357
rect 3141 353 3175 600
rect 3125 319 3175 353
rect 2983 269 3015 319
rect 3143 269 3175 319
rect 2983 217 3017 269
rect 3149 217 3175 269
rect 3183 661 3217 713
rect 3349 679 3375 713
rect 3183 611 3215 661
rect 3325 651 3375 679
rect 3325 645 3341 651
rect 3343 611 3375 651
rect 3183 601 3217 611
rect 3341 601 3375 611
rect 3183 600 3375 601
rect 3183 319 3217 600
rect 3227 573 3251 577
rect 3307 573 3331 577
rect 3221 572 3267 573
rect 3227 353 3251 572
rect 3259 369 3261 561
rect 3263 400 3267 572
rect 3285 572 3337 573
rect 3285 357 3331 572
rect 3307 353 3331 357
rect 3341 353 3375 600
rect 3325 319 3375 353
rect 3183 269 3215 319
rect 3343 269 3375 319
rect 3183 217 3217 269
rect 3349 217 3375 269
rect 3383 661 3417 713
rect 3549 679 3575 713
rect 3383 611 3415 661
rect 3525 651 3575 679
rect 3525 645 3541 651
rect 3543 611 3575 651
rect 3383 601 3417 611
rect 3541 601 3575 611
rect 3383 600 3575 601
rect 3383 319 3417 600
rect 3427 573 3451 577
rect 3507 573 3531 577
rect 3421 572 3467 573
rect 3427 353 3451 572
rect 3459 369 3461 561
rect 3463 400 3467 572
rect 3485 572 3537 573
rect 3485 357 3531 572
rect 3507 353 3531 357
rect 3541 353 3575 600
rect 3525 319 3575 353
rect 3383 269 3415 319
rect 3543 269 3575 319
rect 3383 217 3417 269
rect 3549 217 3575 269
rect 3583 661 3617 713
rect 3583 611 3615 661
rect 3725 651 3775 679
rect 3725 645 3741 651
rect 3743 611 3775 651
rect 3799 611 3809 645
rect 3583 601 3617 611
rect 3741 601 3775 611
rect 3583 600 3775 601
rect 3793 600 3895 601
rect 3583 319 3617 600
rect 3627 573 3651 577
rect 3707 573 3731 577
rect 3621 572 3667 573
rect 3627 353 3651 572
rect 3659 369 3661 561
rect 3663 400 3667 572
rect 3685 572 3737 573
rect 3685 357 3731 572
rect 3707 353 3731 357
rect 3741 353 3775 600
rect 3821 572 3867 573
rect 3725 319 3775 353
rect 3583 269 3615 319
rect 3743 269 3775 319
rect 3799 285 3809 319
rect 3583 217 3617 269
rect 3764 258 3775 269
rect 3947 217 4017 731
rect 4063 600 4165 610
rect 4193 600 4295 610
rect 4091 572 4137 582
rect 4221 572 4267 582
rect 2583 183 2629 217
rect 2679 183 3879 217
rect 3947 183 4029 217
rect 4349 183 4375 749
rect 4383 749 4812 765
rect 4383 731 4429 749
rect 4729 747 4812 749
rect 8947 765 9011 783
rect 9347 765 9412 783
rect 8947 749 9412 765
rect 4383 217 4417 731
rect 4747 713 4829 747
rect 4879 713 6079 747
rect 4463 600 4565 610
rect 4593 600 4695 610
rect 4491 572 4537 582
rect 4621 572 4667 582
rect 4747 217 4817 713
rect 5149 679 5175 713
rect 4983 661 4994 672
rect 4943 611 4959 645
rect 4983 611 5015 661
rect 5125 651 5175 679
rect 5125 645 5141 651
rect 5143 611 5175 651
rect 4983 601 5017 611
rect 5141 601 5175 611
rect 4863 600 4965 601
rect 4983 600 5175 601
rect 4891 572 4937 573
rect 4983 319 5017 600
rect 5027 573 5051 577
rect 5107 573 5131 577
rect 5021 572 5067 573
rect 5027 353 5051 572
rect 5059 369 5061 561
rect 5063 400 5067 572
rect 5085 572 5137 573
rect 5085 357 5131 572
rect 5107 353 5131 357
rect 5141 353 5175 600
rect 5125 319 5175 353
rect 4943 285 4959 319
rect 4983 269 5015 319
rect 5143 269 5175 319
rect 4983 258 4994 269
rect 5149 217 5175 269
rect 5183 661 5217 713
rect 5349 679 5375 713
rect 5183 611 5215 661
rect 5325 651 5375 679
rect 5325 645 5341 651
rect 5343 611 5375 651
rect 5183 601 5217 611
rect 5341 601 5375 611
rect 5183 600 5375 601
rect 5183 319 5217 600
rect 5227 573 5251 577
rect 5307 573 5331 577
rect 5221 572 5267 573
rect 5227 353 5251 572
rect 5259 369 5261 561
rect 5263 400 5267 572
rect 5285 572 5337 573
rect 5285 357 5331 572
rect 5307 353 5331 357
rect 5341 353 5375 600
rect 5325 319 5375 353
rect 5183 269 5215 319
rect 5343 269 5375 319
rect 5183 217 5217 269
rect 5349 217 5375 269
rect 5383 661 5417 713
rect 5549 679 5575 713
rect 5383 611 5415 661
rect 5525 651 5575 679
rect 5525 645 5541 651
rect 5543 611 5575 651
rect 5383 601 5417 611
rect 5541 601 5575 611
rect 5383 600 5575 601
rect 5383 319 5417 600
rect 5427 573 5451 577
rect 5507 573 5531 577
rect 5421 572 5467 573
rect 5427 353 5451 572
rect 5459 369 5461 561
rect 5463 400 5467 572
rect 5485 572 5537 573
rect 5485 357 5531 572
rect 5507 353 5531 357
rect 5541 353 5575 600
rect 5525 319 5575 353
rect 5383 269 5415 319
rect 5543 269 5575 319
rect 5383 217 5417 269
rect 5549 217 5575 269
rect 5583 661 5617 713
rect 5749 679 5775 713
rect 5583 611 5615 661
rect 5725 651 5775 679
rect 5725 645 5741 651
rect 5743 611 5775 651
rect 5583 601 5617 611
rect 5741 601 5775 611
rect 5583 600 5775 601
rect 5583 319 5617 600
rect 5627 573 5651 577
rect 5707 573 5731 577
rect 5621 572 5667 573
rect 5627 353 5651 572
rect 5659 369 5661 561
rect 5663 400 5667 572
rect 5685 572 5737 573
rect 5685 357 5731 572
rect 5707 353 5731 357
rect 5741 353 5775 600
rect 5725 319 5775 353
rect 5583 269 5615 319
rect 5743 269 5775 319
rect 5583 217 5617 269
rect 5749 217 5775 269
rect 5783 661 5817 713
rect 5783 611 5815 661
rect 5925 651 5975 679
rect 5925 645 5941 651
rect 5943 611 5975 651
rect 5999 611 6009 645
rect 5783 601 5817 611
rect 5941 601 5975 611
rect 5783 600 5975 601
rect 5993 600 6095 601
rect 5783 319 5817 600
rect 5827 573 5851 577
rect 5907 573 5931 577
rect 5821 572 5867 573
rect 5827 353 5851 572
rect 5859 369 5861 561
rect 5863 400 5867 572
rect 5885 572 5937 573
rect 5885 357 5931 572
rect 5907 353 5931 357
rect 5941 353 5975 600
rect 6021 572 6067 573
rect 5925 319 5975 353
rect 5783 269 5815 319
rect 5943 269 5975 319
rect 5999 285 6009 319
rect 5783 217 5817 269
rect 5964 258 5975 269
rect 4383 183 4429 217
rect 4747 183 4829 217
rect 4879 183 6079 217
rect 6149 183 6175 747
rect 6183 713 6229 747
rect 6279 713 7479 747
rect 6183 217 6217 713
rect 6549 679 6575 713
rect 6383 661 6394 672
rect 6343 611 6359 645
rect 6383 611 6415 661
rect 6525 651 6575 679
rect 6525 645 6541 651
rect 6543 611 6575 651
rect 6383 601 6417 611
rect 6541 601 6575 611
rect 6263 600 6365 601
rect 6383 600 6575 601
rect 6291 572 6337 573
rect 6383 319 6417 600
rect 6427 573 6451 577
rect 6507 573 6531 577
rect 6421 572 6467 573
rect 6427 353 6451 572
rect 6459 369 6461 561
rect 6463 400 6467 572
rect 6485 572 6537 573
rect 6485 357 6531 572
rect 6507 353 6531 357
rect 6541 353 6575 600
rect 6525 319 6575 353
rect 6343 285 6359 319
rect 6383 269 6415 319
rect 6543 269 6575 319
rect 6383 258 6394 269
rect 6549 217 6575 269
rect 6583 661 6617 713
rect 6749 679 6775 713
rect 6583 611 6615 661
rect 6725 651 6775 679
rect 6725 645 6741 651
rect 6743 611 6775 651
rect 6583 601 6617 611
rect 6741 601 6775 611
rect 6583 600 6775 601
rect 6583 319 6617 600
rect 6627 573 6651 577
rect 6707 573 6731 577
rect 6621 572 6667 573
rect 6627 353 6651 572
rect 6659 369 6661 561
rect 6663 400 6667 572
rect 6685 572 6737 573
rect 6685 357 6731 572
rect 6707 353 6731 357
rect 6741 353 6775 600
rect 6725 319 6775 353
rect 6583 269 6615 319
rect 6743 269 6775 319
rect 6583 217 6617 269
rect 6749 217 6775 269
rect 6783 661 6817 713
rect 6949 679 6975 713
rect 6783 611 6815 661
rect 6925 651 6975 679
rect 6925 645 6941 651
rect 6943 611 6975 651
rect 6783 601 6817 611
rect 6941 601 6975 611
rect 6783 600 6975 601
rect 6783 319 6817 600
rect 6827 573 6851 577
rect 6907 573 6931 577
rect 6821 572 6867 573
rect 6827 353 6851 572
rect 6859 369 6861 561
rect 6863 400 6867 572
rect 6885 572 6937 573
rect 6885 357 6931 572
rect 6907 353 6931 357
rect 6941 353 6975 600
rect 6925 319 6975 353
rect 6783 269 6815 319
rect 6943 269 6975 319
rect 6783 217 6817 269
rect 6949 217 6975 269
rect 6983 661 7017 713
rect 7149 679 7175 713
rect 6983 611 7015 661
rect 7125 651 7175 679
rect 7125 645 7141 651
rect 7143 611 7175 651
rect 6983 601 7017 611
rect 7141 601 7175 611
rect 6983 600 7175 601
rect 6983 319 7017 600
rect 7027 573 7051 577
rect 7107 573 7131 577
rect 7021 572 7067 573
rect 7027 353 7051 572
rect 7059 369 7061 561
rect 7063 400 7067 572
rect 7085 572 7137 573
rect 7085 357 7131 572
rect 7107 353 7131 357
rect 7141 353 7175 600
rect 7125 319 7175 353
rect 6983 269 7015 319
rect 7143 269 7175 319
rect 6983 217 7017 269
rect 7149 217 7175 269
rect 7183 661 7217 713
rect 7183 611 7215 661
rect 7325 651 7375 679
rect 7325 645 7341 651
rect 7343 611 7375 651
rect 7399 611 7409 645
rect 7183 601 7217 611
rect 7341 601 7375 611
rect 7183 600 7375 601
rect 7393 600 7495 601
rect 7183 319 7217 600
rect 7227 573 7251 577
rect 7307 573 7331 577
rect 7221 572 7267 573
rect 7227 353 7251 572
rect 7259 369 7261 561
rect 7263 400 7267 572
rect 7285 572 7337 573
rect 7285 357 7331 572
rect 7307 353 7331 357
rect 7341 353 7375 600
rect 7421 572 7467 573
rect 7325 319 7375 353
rect 7183 269 7215 319
rect 7343 269 7375 319
rect 7399 285 7409 319
rect 7183 217 7217 269
rect 7364 258 7375 269
rect 6183 183 6229 217
rect 6279 183 7479 217
rect 7549 183 7575 747
rect 7583 713 7629 747
rect 7679 713 8879 747
rect 8947 731 9029 749
rect 9329 747 9412 749
rect 10747 765 10811 783
rect 11147 765 11212 783
rect 10747 749 11212 765
rect 7583 217 7617 713
rect 7949 679 7975 713
rect 7783 661 7794 672
rect 7743 611 7759 645
rect 7783 611 7815 661
rect 7925 651 7975 679
rect 7925 645 7941 651
rect 7943 611 7975 651
rect 7783 601 7817 611
rect 7941 601 7975 611
rect 7663 600 7765 601
rect 7783 600 7975 601
rect 7691 572 7737 573
rect 7783 319 7817 600
rect 7827 573 7851 577
rect 7907 573 7931 577
rect 7821 572 7867 573
rect 7827 353 7851 572
rect 7859 369 7861 561
rect 7863 400 7867 572
rect 7885 572 7937 573
rect 7885 357 7931 572
rect 7907 353 7931 357
rect 7941 353 7975 600
rect 7925 319 7975 353
rect 7743 285 7759 319
rect 7783 269 7815 319
rect 7943 269 7975 319
rect 7783 258 7794 269
rect 7949 217 7975 269
rect 7983 661 8017 713
rect 8149 679 8175 713
rect 7983 611 8015 661
rect 8125 651 8175 679
rect 8125 645 8141 651
rect 8143 611 8175 651
rect 7983 601 8017 611
rect 8141 601 8175 611
rect 7983 600 8175 601
rect 7983 319 8017 600
rect 8027 573 8051 577
rect 8107 573 8131 577
rect 8021 572 8067 573
rect 8027 353 8051 572
rect 8059 369 8061 561
rect 8063 400 8067 572
rect 8085 572 8137 573
rect 8085 357 8131 572
rect 8107 353 8131 357
rect 8141 353 8175 600
rect 8125 319 8175 353
rect 7983 269 8015 319
rect 8143 269 8175 319
rect 7983 217 8017 269
rect 8149 217 8175 269
rect 8183 661 8217 713
rect 8349 679 8375 713
rect 8183 611 8215 661
rect 8325 651 8375 679
rect 8325 645 8341 651
rect 8343 611 8375 651
rect 8183 601 8217 611
rect 8341 601 8375 611
rect 8183 600 8375 601
rect 8183 319 8217 600
rect 8227 573 8251 577
rect 8307 573 8331 577
rect 8221 572 8267 573
rect 8227 353 8251 572
rect 8259 369 8261 561
rect 8263 400 8267 572
rect 8285 572 8337 573
rect 8285 357 8331 572
rect 8307 353 8331 357
rect 8341 353 8375 600
rect 8325 319 8375 353
rect 8183 269 8215 319
rect 8343 269 8375 319
rect 8183 217 8217 269
rect 8349 217 8375 269
rect 8383 661 8417 713
rect 8549 679 8575 713
rect 8383 611 8415 661
rect 8525 651 8575 679
rect 8525 645 8541 651
rect 8543 611 8575 651
rect 8383 601 8417 611
rect 8541 601 8575 611
rect 8383 600 8575 601
rect 8383 319 8417 600
rect 8427 573 8451 577
rect 8507 573 8531 577
rect 8421 572 8467 573
rect 8427 353 8451 572
rect 8459 369 8461 561
rect 8463 400 8467 572
rect 8485 572 8537 573
rect 8485 357 8531 572
rect 8507 353 8531 357
rect 8541 353 8575 600
rect 8525 319 8575 353
rect 8383 269 8415 319
rect 8543 269 8575 319
rect 8383 217 8417 269
rect 8549 217 8575 269
rect 8583 661 8617 713
rect 8583 611 8615 661
rect 8725 651 8775 679
rect 8725 645 8741 651
rect 8743 611 8775 651
rect 8799 611 8809 645
rect 8583 601 8617 611
rect 8741 601 8775 611
rect 8583 600 8775 601
rect 8793 600 8895 601
rect 8583 319 8617 600
rect 8627 573 8651 577
rect 8707 573 8731 577
rect 8621 572 8667 573
rect 8627 353 8651 572
rect 8659 369 8661 561
rect 8663 400 8667 572
rect 8685 572 8737 573
rect 8685 357 8731 572
rect 8707 353 8731 357
rect 8741 353 8775 600
rect 8821 572 8867 573
rect 8725 319 8775 353
rect 8583 269 8615 319
rect 8743 269 8775 319
rect 8799 285 8809 319
rect 8583 217 8617 269
rect 8764 258 8775 269
rect 8947 217 9017 731
rect 9347 713 9429 747
rect 9479 713 10679 747
rect 10747 731 10829 749
rect 11129 747 11212 749
rect 12547 765 12611 783
rect 12947 765 13012 783
rect 12547 749 13012 765
rect 9063 600 9165 610
rect 9193 600 9295 610
rect 9091 572 9137 582
rect 9221 572 9267 582
rect 9347 217 9417 713
rect 9749 679 9775 713
rect 9583 661 9594 672
rect 9543 611 9559 645
rect 9583 611 9615 661
rect 9725 651 9775 679
rect 9725 645 9741 651
rect 9743 611 9775 651
rect 9583 601 9617 611
rect 9741 601 9775 611
rect 9463 600 9565 601
rect 9583 600 9775 601
rect 9491 572 9537 573
rect 9583 319 9617 600
rect 9627 573 9651 577
rect 9707 573 9731 577
rect 9621 572 9667 573
rect 9627 353 9651 572
rect 9659 369 9661 561
rect 9663 400 9667 572
rect 9685 572 9737 573
rect 9685 357 9731 572
rect 9707 353 9731 357
rect 9741 353 9775 600
rect 9725 319 9775 353
rect 9543 285 9559 319
rect 9583 269 9615 319
rect 9743 269 9775 319
rect 9583 258 9594 269
rect 9749 217 9775 269
rect 9783 661 9817 713
rect 9949 679 9975 713
rect 9783 611 9815 661
rect 9925 651 9975 679
rect 9925 645 9941 651
rect 9943 611 9975 651
rect 9783 601 9817 611
rect 9941 601 9975 611
rect 9783 600 9975 601
rect 9783 319 9817 600
rect 9827 573 9851 577
rect 9907 573 9931 577
rect 9821 572 9867 573
rect 9827 353 9851 572
rect 9859 369 9861 561
rect 9863 400 9867 572
rect 9885 572 9937 573
rect 9885 357 9931 572
rect 9907 353 9931 357
rect 9941 353 9975 600
rect 9925 319 9975 353
rect 9783 269 9815 319
rect 9943 269 9975 319
rect 9783 217 9817 269
rect 9949 217 9975 269
rect 9983 661 10017 713
rect 10149 679 10175 713
rect 9983 611 10015 661
rect 10125 651 10175 679
rect 10125 645 10141 651
rect 10143 611 10175 651
rect 9983 601 10017 611
rect 10141 601 10175 611
rect 9983 600 10175 601
rect 9983 319 10017 600
rect 10027 573 10051 577
rect 10107 573 10131 577
rect 10021 572 10067 573
rect 10027 353 10051 572
rect 10059 369 10061 561
rect 10063 400 10067 572
rect 10085 572 10137 573
rect 10085 357 10131 572
rect 10107 353 10131 357
rect 10141 353 10175 600
rect 10125 319 10175 353
rect 9983 269 10015 319
rect 10143 269 10175 319
rect 9983 217 10017 269
rect 10149 217 10175 269
rect 10183 661 10217 713
rect 10349 679 10375 713
rect 10183 611 10215 661
rect 10325 651 10375 679
rect 10325 645 10341 651
rect 10343 611 10375 651
rect 10183 601 10217 611
rect 10341 601 10375 611
rect 10183 600 10375 601
rect 10183 319 10217 600
rect 10227 573 10251 577
rect 10307 573 10331 577
rect 10221 572 10267 573
rect 10227 353 10251 572
rect 10259 369 10261 561
rect 10263 400 10267 572
rect 10285 572 10337 573
rect 10285 357 10331 572
rect 10307 353 10331 357
rect 10341 353 10375 600
rect 10325 319 10375 353
rect 10183 269 10215 319
rect 10343 269 10375 319
rect 10183 217 10217 269
rect 10349 217 10375 269
rect 10383 661 10417 713
rect 10383 611 10415 661
rect 10525 651 10575 679
rect 10525 645 10541 651
rect 10543 611 10575 651
rect 10599 611 10609 645
rect 10383 601 10417 611
rect 10541 601 10575 611
rect 10383 600 10575 601
rect 10593 600 10695 601
rect 10383 319 10417 600
rect 10427 573 10451 577
rect 10507 573 10531 577
rect 10421 572 10467 573
rect 10427 353 10451 572
rect 10459 369 10461 561
rect 10463 400 10467 572
rect 10485 572 10537 573
rect 10485 357 10531 572
rect 10507 353 10531 357
rect 10541 353 10575 600
rect 10621 572 10667 573
rect 10525 319 10575 353
rect 10383 269 10415 319
rect 10543 269 10575 319
rect 10599 285 10609 319
rect 10383 217 10417 269
rect 10564 258 10575 269
rect 10747 217 10817 731
rect 11147 713 11229 747
rect 11279 713 12479 747
rect 12547 731 12629 749
rect 12929 747 13012 749
rect 14347 765 14411 783
rect 14747 765 14812 783
rect 14347 749 14812 765
rect 10863 600 10965 610
rect 10993 600 11095 610
rect 10891 572 10937 582
rect 11021 572 11067 582
rect 11147 217 11217 713
rect 11549 679 11575 713
rect 11383 661 11394 672
rect 11343 611 11359 645
rect 11383 611 11415 661
rect 11525 651 11575 679
rect 11525 645 11541 651
rect 11543 611 11575 651
rect 11383 601 11417 611
rect 11541 601 11575 611
rect 11263 600 11365 601
rect 11383 600 11575 601
rect 11291 572 11337 573
rect 11383 319 11417 600
rect 11427 573 11451 577
rect 11507 573 11531 577
rect 11421 572 11467 573
rect 11427 353 11451 572
rect 11459 369 11461 561
rect 11463 400 11467 572
rect 11485 572 11537 573
rect 11485 357 11531 572
rect 11507 353 11531 357
rect 11541 353 11575 600
rect 11525 319 11575 353
rect 11343 285 11359 319
rect 11383 269 11415 319
rect 11543 269 11575 319
rect 11383 258 11394 269
rect 11549 217 11575 269
rect 11583 661 11617 713
rect 11749 679 11775 713
rect 11583 611 11615 661
rect 11725 651 11775 679
rect 11725 645 11741 651
rect 11743 611 11775 651
rect 11583 601 11617 611
rect 11741 601 11775 611
rect 11583 600 11775 601
rect 11583 319 11617 600
rect 11627 573 11651 577
rect 11707 573 11731 577
rect 11621 572 11667 573
rect 11627 353 11651 572
rect 11659 369 11661 561
rect 11663 400 11667 572
rect 11685 572 11737 573
rect 11685 357 11731 572
rect 11707 353 11731 357
rect 11741 353 11775 600
rect 11725 319 11775 353
rect 11583 269 11615 319
rect 11743 269 11775 319
rect 11583 217 11617 269
rect 11749 217 11775 269
rect 11783 661 11817 713
rect 11949 679 11975 713
rect 11783 611 11815 661
rect 11925 651 11975 679
rect 11925 645 11941 651
rect 11943 611 11975 651
rect 11783 601 11817 611
rect 11941 601 11975 611
rect 11783 600 11975 601
rect 11783 319 11817 600
rect 11827 573 11851 577
rect 11907 573 11931 577
rect 11821 572 11867 573
rect 11827 353 11851 572
rect 11859 369 11861 561
rect 11863 400 11867 572
rect 11885 572 11937 573
rect 11885 357 11931 572
rect 11907 353 11931 357
rect 11941 353 11975 600
rect 11925 319 11975 353
rect 11783 269 11815 319
rect 11943 269 11975 319
rect 11783 217 11817 269
rect 11949 217 11975 269
rect 11983 661 12017 713
rect 12149 679 12175 713
rect 11983 611 12015 661
rect 12125 651 12175 679
rect 12125 645 12141 651
rect 12143 611 12175 651
rect 11983 601 12017 611
rect 12141 601 12175 611
rect 11983 600 12175 601
rect 11983 319 12017 600
rect 12027 573 12051 577
rect 12107 573 12131 577
rect 12021 572 12067 573
rect 12027 353 12051 572
rect 12059 369 12061 561
rect 12063 400 12067 572
rect 12085 572 12137 573
rect 12085 357 12131 572
rect 12107 353 12131 357
rect 12141 353 12175 600
rect 12125 319 12175 353
rect 11983 269 12015 319
rect 12143 269 12175 319
rect 11983 217 12017 269
rect 12149 217 12175 269
rect 12183 661 12217 713
rect 12183 611 12215 661
rect 12325 651 12375 679
rect 12325 645 12341 651
rect 12343 611 12375 651
rect 12399 611 12409 645
rect 12183 601 12217 611
rect 12341 601 12375 611
rect 12183 600 12375 601
rect 12393 600 12495 601
rect 12183 319 12217 600
rect 12227 573 12251 577
rect 12307 573 12331 577
rect 12221 572 12267 573
rect 12227 353 12251 572
rect 12259 369 12261 561
rect 12263 400 12267 572
rect 12285 572 12337 573
rect 12285 357 12331 572
rect 12307 353 12331 357
rect 12341 353 12375 600
rect 12421 572 12467 573
rect 12325 319 12375 353
rect 12183 269 12215 319
rect 12343 269 12375 319
rect 12399 285 12409 319
rect 12183 217 12217 269
rect 12364 258 12375 269
rect 12547 217 12617 731
rect 12947 713 13029 747
rect 13079 713 14279 747
rect 14347 731 14429 749
rect 14729 747 14812 749
rect 16147 765 16211 783
rect 16547 765 16612 783
rect 16147 749 16612 765
rect 12663 600 12765 610
rect 12793 600 12895 610
rect 12691 572 12737 582
rect 12821 572 12867 582
rect 12947 217 13017 713
rect 13349 679 13375 713
rect 13183 661 13194 672
rect 13143 611 13159 645
rect 13183 611 13215 661
rect 13325 651 13375 679
rect 13325 645 13341 651
rect 13343 611 13375 651
rect 13183 601 13217 611
rect 13341 601 13375 611
rect 13063 600 13165 601
rect 13183 600 13375 601
rect 13091 572 13137 573
rect 13183 319 13217 600
rect 13227 573 13251 577
rect 13307 573 13331 577
rect 13221 572 13267 573
rect 13227 353 13251 572
rect 13259 369 13261 561
rect 13263 400 13267 572
rect 13285 572 13337 573
rect 13285 357 13331 572
rect 13307 353 13331 357
rect 13341 353 13375 600
rect 13325 319 13375 353
rect 13143 285 13159 319
rect 13183 269 13215 319
rect 13343 269 13375 319
rect 13183 258 13194 269
rect 13349 217 13375 269
rect 13383 661 13417 713
rect 13549 679 13575 713
rect 13383 611 13415 661
rect 13525 651 13575 679
rect 13525 645 13541 651
rect 13543 611 13575 651
rect 13383 601 13417 611
rect 13541 601 13575 611
rect 13383 600 13575 601
rect 13383 319 13417 600
rect 13427 573 13451 577
rect 13507 573 13531 577
rect 13421 572 13467 573
rect 13427 353 13451 572
rect 13459 369 13461 561
rect 13463 400 13467 572
rect 13485 572 13537 573
rect 13485 357 13531 572
rect 13507 353 13531 357
rect 13541 353 13575 600
rect 13525 319 13575 353
rect 13383 269 13415 319
rect 13543 269 13575 319
rect 13383 217 13417 269
rect 13549 217 13575 269
rect 13583 661 13617 713
rect 13749 679 13775 713
rect 13583 611 13615 661
rect 13725 651 13775 679
rect 13725 645 13741 651
rect 13743 611 13775 651
rect 13583 601 13617 611
rect 13741 601 13775 611
rect 13583 600 13775 601
rect 13583 319 13617 600
rect 13627 573 13651 577
rect 13707 573 13731 577
rect 13621 572 13667 573
rect 13627 353 13651 572
rect 13659 369 13661 561
rect 13663 400 13667 572
rect 13685 572 13737 573
rect 13685 357 13731 572
rect 13707 353 13731 357
rect 13741 353 13775 600
rect 13725 319 13775 353
rect 13583 269 13615 319
rect 13743 269 13775 319
rect 13583 217 13617 269
rect 13749 217 13775 269
rect 13783 661 13817 713
rect 13949 679 13975 713
rect 13783 611 13815 661
rect 13925 651 13975 679
rect 13925 645 13941 651
rect 13943 611 13975 651
rect 13783 601 13817 611
rect 13941 601 13975 611
rect 13783 600 13975 601
rect 13783 319 13817 600
rect 13827 573 13851 577
rect 13907 573 13931 577
rect 13821 572 13867 573
rect 13827 353 13851 572
rect 13859 369 13861 561
rect 13863 400 13867 572
rect 13885 572 13937 573
rect 13885 357 13931 572
rect 13907 353 13931 357
rect 13941 353 13975 600
rect 13925 319 13975 353
rect 13783 269 13815 319
rect 13943 269 13975 319
rect 13783 217 13817 269
rect 13949 217 13975 269
rect 13983 661 14017 713
rect 13983 611 14015 661
rect 14125 651 14175 679
rect 14125 645 14141 651
rect 14143 611 14175 651
rect 14199 611 14209 645
rect 13983 601 14017 611
rect 14141 601 14175 611
rect 13983 600 14175 601
rect 14193 600 14295 601
rect 13983 319 14017 600
rect 14027 573 14051 577
rect 14107 573 14131 577
rect 14021 572 14067 573
rect 14027 353 14051 572
rect 14059 369 14061 561
rect 14063 400 14067 572
rect 14085 572 14137 573
rect 14085 357 14131 572
rect 14107 353 14131 357
rect 14141 353 14175 600
rect 14221 572 14267 573
rect 14125 319 14175 353
rect 13983 269 14015 319
rect 14143 269 14175 319
rect 14199 285 14209 319
rect 13983 217 14017 269
rect 14164 258 14175 269
rect 14347 217 14417 731
rect 14747 713 14829 747
rect 14879 713 16079 747
rect 16147 731 16229 749
rect 16529 747 16612 749
rect 19347 765 19411 783
rect 20147 765 20212 783
rect 19347 749 19775 765
rect 14463 600 14565 610
rect 14593 600 14695 610
rect 14491 572 14537 582
rect 14621 572 14667 582
rect 14747 217 14817 713
rect 15149 679 15175 713
rect 14983 661 14994 672
rect 14943 611 14959 645
rect 14983 611 15015 661
rect 15125 651 15175 679
rect 15125 645 15141 651
rect 15143 611 15175 651
rect 14983 601 15017 611
rect 15141 601 15175 611
rect 14863 600 14965 601
rect 14983 600 15175 601
rect 14891 572 14937 573
rect 14983 319 15017 600
rect 15027 573 15051 577
rect 15107 573 15131 577
rect 15021 572 15067 573
rect 15027 353 15051 572
rect 15059 369 15061 561
rect 15063 400 15067 572
rect 15085 572 15137 573
rect 15085 357 15131 572
rect 15107 353 15131 357
rect 15141 353 15175 600
rect 15125 319 15175 353
rect 14943 285 14959 319
rect 14983 269 15015 319
rect 15143 269 15175 319
rect 14983 258 14994 269
rect 15149 217 15175 269
rect 15183 661 15217 713
rect 15349 679 15375 713
rect 15183 611 15215 661
rect 15325 651 15375 679
rect 15325 645 15341 651
rect 15343 611 15375 651
rect 15183 601 15217 611
rect 15341 601 15375 611
rect 15183 600 15375 601
rect 15183 319 15217 600
rect 15227 573 15251 577
rect 15307 573 15331 577
rect 15221 572 15267 573
rect 15227 353 15251 572
rect 15259 369 15261 561
rect 15263 400 15267 572
rect 15285 572 15337 573
rect 15285 357 15331 572
rect 15307 353 15331 357
rect 15341 353 15375 600
rect 15325 319 15375 353
rect 15183 269 15215 319
rect 15343 269 15375 319
rect 15183 217 15217 269
rect 15349 217 15375 269
rect 15383 661 15417 713
rect 15549 679 15575 713
rect 15383 611 15415 661
rect 15525 651 15575 679
rect 15525 645 15541 651
rect 15543 611 15575 651
rect 15383 601 15417 611
rect 15541 601 15575 611
rect 15383 600 15575 601
rect 15383 319 15417 600
rect 15427 573 15451 577
rect 15507 573 15531 577
rect 15421 572 15467 573
rect 15427 353 15451 572
rect 15459 369 15461 561
rect 15463 400 15467 572
rect 15485 572 15537 573
rect 15485 357 15531 572
rect 15507 353 15531 357
rect 15541 353 15575 600
rect 15525 319 15575 353
rect 15383 269 15415 319
rect 15543 269 15575 319
rect 15383 217 15417 269
rect 15549 217 15575 269
rect 15583 661 15617 713
rect 15749 679 15775 713
rect 15583 611 15615 661
rect 15725 651 15775 679
rect 15725 645 15741 651
rect 15743 611 15775 651
rect 15583 601 15617 611
rect 15741 601 15775 611
rect 15583 600 15775 601
rect 15583 319 15617 600
rect 15627 573 15651 577
rect 15707 573 15731 577
rect 15621 572 15667 573
rect 15627 353 15651 572
rect 15659 369 15661 561
rect 15663 400 15667 572
rect 15685 572 15737 573
rect 15685 357 15731 572
rect 15707 353 15731 357
rect 15741 353 15775 600
rect 15725 319 15775 353
rect 15583 269 15615 319
rect 15743 269 15775 319
rect 15583 217 15617 269
rect 15749 217 15775 269
rect 15783 661 15817 713
rect 15783 611 15815 661
rect 15925 651 15975 679
rect 15925 645 15941 651
rect 15943 611 15975 651
rect 15999 611 16009 645
rect 15783 601 15817 611
rect 15941 601 15975 611
rect 15783 600 15975 601
rect 15993 600 16095 601
rect 15783 319 15817 600
rect 15827 573 15851 577
rect 15907 573 15931 577
rect 15821 572 15867 573
rect 15827 353 15851 572
rect 15859 369 15861 561
rect 15863 400 15867 572
rect 15885 572 15937 573
rect 15885 357 15931 572
rect 15907 353 15931 357
rect 15941 353 15975 600
rect 16021 572 16067 573
rect 15925 319 15975 353
rect 15783 269 15815 319
rect 15943 269 15975 319
rect 15999 285 16009 319
rect 15783 217 15817 269
rect 15964 258 15975 269
rect 16147 217 16217 731
rect 16547 713 16629 747
rect 16679 713 17879 747
rect 16263 600 16365 610
rect 16393 600 16495 610
rect 16291 572 16337 582
rect 16421 572 16467 582
rect 16547 217 16617 713
rect 16949 679 16975 713
rect 16783 661 16794 672
rect 16743 611 16759 645
rect 16783 611 16815 661
rect 16925 651 16975 679
rect 16925 645 16941 651
rect 16943 611 16975 651
rect 16783 601 16817 611
rect 16941 601 16975 611
rect 16663 600 16765 601
rect 16783 600 16975 601
rect 16691 572 16737 573
rect 16783 319 16817 600
rect 16827 573 16851 577
rect 16907 573 16931 577
rect 16821 572 16867 573
rect 16827 353 16851 572
rect 16859 369 16861 561
rect 16863 400 16867 572
rect 16885 572 16937 573
rect 16885 357 16931 572
rect 16907 353 16931 357
rect 16941 353 16975 600
rect 16925 319 16975 353
rect 16743 285 16759 319
rect 16783 269 16815 319
rect 16943 269 16975 319
rect 16783 258 16794 269
rect 16949 217 16975 269
rect 16983 661 17017 713
rect 17149 679 17175 713
rect 16983 611 17015 661
rect 17125 651 17175 679
rect 17125 645 17141 651
rect 17143 611 17175 651
rect 16983 601 17017 611
rect 17141 601 17175 611
rect 16983 600 17175 601
rect 16983 319 17017 600
rect 17027 573 17051 577
rect 17107 573 17131 577
rect 17021 572 17067 573
rect 17027 353 17051 572
rect 17059 369 17061 561
rect 17063 400 17067 572
rect 17085 572 17137 573
rect 17085 357 17131 572
rect 17107 353 17131 357
rect 17141 353 17175 600
rect 17125 319 17175 353
rect 16983 269 17015 319
rect 17143 269 17175 319
rect 16983 217 17017 269
rect 17149 217 17175 269
rect 17183 661 17217 713
rect 17349 679 17375 713
rect 17183 611 17215 661
rect 17325 651 17375 679
rect 17325 645 17341 651
rect 17343 611 17375 651
rect 17183 601 17217 611
rect 17341 601 17375 611
rect 17183 600 17375 601
rect 17183 319 17217 600
rect 17227 573 17251 577
rect 17307 573 17331 577
rect 17221 572 17267 573
rect 17227 353 17251 572
rect 17259 369 17261 561
rect 17263 400 17267 572
rect 17285 572 17337 573
rect 17285 357 17331 572
rect 17307 353 17331 357
rect 17341 353 17375 600
rect 17325 319 17375 353
rect 17183 269 17215 319
rect 17343 269 17375 319
rect 17183 217 17217 269
rect 17349 217 17375 269
rect 17383 661 17417 713
rect 17549 679 17575 713
rect 17383 611 17415 661
rect 17525 651 17575 679
rect 17525 645 17541 651
rect 17543 611 17575 651
rect 17383 601 17417 611
rect 17541 601 17575 611
rect 17383 600 17575 601
rect 17383 319 17417 600
rect 17427 573 17451 577
rect 17507 573 17531 577
rect 17421 572 17467 573
rect 17427 353 17451 572
rect 17459 369 17461 561
rect 17463 400 17467 572
rect 17485 572 17537 573
rect 17485 357 17531 572
rect 17507 353 17531 357
rect 17541 353 17575 600
rect 17525 319 17575 353
rect 17383 269 17415 319
rect 17543 269 17575 319
rect 17383 217 17417 269
rect 17549 217 17575 269
rect 17583 661 17617 713
rect 17583 611 17615 661
rect 17725 651 17775 679
rect 17725 645 17741 651
rect 17743 611 17775 651
rect 17799 611 17809 645
rect 17583 601 17617 611
rect 17741 601 17775 611
rect 17583 600 17775 601
rect 17793 600 17895 601
rect 17583 319 17617 600
rect 17627 573 17651 577
rect 17707 573 17731 577
rect 17621 572 17667 573
rect 17627 353 17651 572
rect 17659 369 17661 561
rect 17663 400 17667 572
rect 17685 572 17737 573
rect 17685 357 17731 572
rect 17707 353 17731 357
rect 17741 353 17775 600
rect 17821 572 17867 573
rect 17725 319 17775 353
rect 17583 269 17615 319
rect 17743 269 17775 319
rect 17799 285 17809 319
rect 17583 217 17617 269
rect 17764 258 17775 269
rect 7583 183 7629 217
rect 7679 183 8879 217
rect 8947 183 9029 217
rect 9347 183 9429 217
rect 9479 183 10679 217
rect 10747 183 10829 217
rect 11147 183 11229 217
rect 11279 183 12479 217
rect 12547 183 12629 217
rect 12947 183 13029 217
rect 13079 183 14279 217
rect 14347 183 14429 217
rect 14747 183 14829 217
rect 14879 183 16079 217
rect 16147 183 16229 217
rect 16547 183 16629 217
rect 16679 183 17879 217
rect 17949 183 17975 747
rect 17983 713 18029 747
rect 18079 713 19279 747
rect 19347 731 19429 749
rect 17983 217 18017 713
rect 18349 679 18375 713
rect 18183 661 18194 672
rect 18143 611 18159 645
rect 18183 611 18215 661
rect 18325 651 18375 679
rect 18325 645 18341 651
rect 18343 611 18375 651
rect 18183 601 18217 611
rect 18341 601 18375 611
rect 18063 600 18165 601
rect 18183 600 18375 601
rect 18091 572 18137 573
rect 18183 319 18217 600
rect 18227 573 18251 577
rect 18307 573 18331 577
rect 18221 572 18267 573
rect 18227 353 18251 572
rect 18259 369 18261 561
rect 18263 400 18267 572
rect 18285 572 18337 573
rect 18285 357 18331 572
rect 18307 353 18331 357
rect 18341 353 18375 600
rect 18325 319 18375 353
rect 18143 285 18159 319
rect 18183 269 18215 319
rect 18343 269 18375 319
rect 18183 258 18194 269
rect 18349 217 18375 269
rect 18383 661 18417 713
rect 18549 679 18575 713
rect 18383 611 18415 661
rect 18525 651 18575 679
rect 18525 645 18541 651
rect 18543 611 18575 651
rect 18383 601 18417 611
rect 18541 601 18575 611
rect 18383 600 18575 601
rect 18383 319 18417 600
rect 18427 573 18451 577
rect 18507 573 18531 577
rect 18421 572 18467 573
rect 18427 353 18451 572
rect 18459 369 18461 561
rect 18463 400 18467 572
rect 18485 572 18537 573
rect 18485 357 18531 572
rect 18507 353 18531 357
rect 18541 353 18575 600
rect 18525 319 18575 353
rect 18383 269 18415 319
rect 18543 269 18575 319
rect 18383 217 18417 269
rect 18549 217 18575 269
rect 18583 661 18617 713
rect 18749 679 18775 713
rect 18583 611 18615 661
rect 18725 651 18775 679
rect 18725 645 18741 651
rect 18743 611 18775 651
rect 18583 601 18617 611
rect 18741 601 18775 611
rect 18583 600 18775 601
rect 18583 319 18617 600
rect 18627 573 18651 577
rect 18707 573 18731 577
rect 18621 572 18667 573
rect 18627 353 18651 572
rect 18659 369 18661 561
rect 18663 400 18667 572
rect 18685 572 18737 573
rect 18685 357 18731 572
rect 18707 353 18731 357
rect 18741 353 18775 600
rect 18725 319 18775 353
rect 18583 269 18615 319
rect 18743 269 18775 319
rect 18583 217 18617 269
rect 18749 217 18775 269
rect 18783 661 18817 713
rect 18949 679 18975 713
rect 18783 611 18815 661
rect 18925 651 18975 679
rect 18925 645 18941 651
rect 18943 611 18975 651
rect 18783 601 18817 611
rect 18941 601 18975 611
rect 18783 600 18975 601
rect 18783 319 18817 600
rect 18827 573 18851 577
rect 18907 573 18931 577
rect 18821 572 18867 573
rect 18827 353 18851 572
rect 18859 369 18861 561
rect 18863 400 18867 572
rect 18885 572 18937 573
rect 18885 357 18931 572
rect 18907 353 18931 357
rect 18941 353 18975 600
rect 18925 319 18975 353
rect 18783 269 18815 319
rect 18943 269 18975 319
rect 18783 217 18817 269
rect 18949 217 18975 269
rect 18983 661 19017 713
rect 18983 611 19015 661
rect 19125 651 19175 679
rect 19125 645 19141 651
rect 19143 611 19175 651
rect 19199 611 19209 645
rect 18983 601 19017 611
rect 19141 601 19175 611
rect 18983 600 19175 601
rect 19193 600 19295 601
rect 18983 319 19017 600
rect 19027 573 19051 577
rect 19107 573 19131 577
rect 19021 572 19067 573
rect 19027 353 19051 572
rect 19059 369 19061 561
rect 19063 400 19067 572
rect 19085 572 19137 573
rect 19085 357 19131 572
rect 19107 353 19131 357
rect 19141 353 19175 600
rect 19221 572 19267 573
rect 19125 319 19175 353
rect 18983 269 19015 319
rect 19143 269 19175 319
rect 19199 285 19209 319
rect 18983 217 19017 269
rect 19164 258 19175 269
rect 19347 217 19417 731
rect 19463 600 19565 610
rect 19593 600 19695 610
rect 19491 572 19537 582
rect 19621 572 19667 582
rect 17983 183 18029 217
rect 18079 183 19279 217
rect 19347 183 19429 217
rect 19749 183 19775 749
rect 19783 749 20212 765
rect 19783 731 19829 749
rect 20129 747 20212 749
rect 21547 765 21611 783
rect 21947 765 22012 783
rect 21547 749 22012 765
rect 19783 217 19817 731
rect 20147 713 20229 747
rect 20279 713 21479 747
rect 21547 731 21629 749
rect 21929 747 22012 749
rect 23347 765 23411 783
rect 23747 765 23812 783
rect 23347 749 23812 765
rect 19863 600 19965 610
rect 19993 600 20095 610
rect 19891 572 19937 582
rect 20021 572 20067 582
rect 20147 217 20217 713
rect 20549 679 20575 713
rect 20383 661 20394 672
rect 20343 611 20359 645
rect 20383 611 20415 661
rect 20525 651 20575 679
rect 20525 645 20541 651
rect 20543 611 20575 651
rect 20383 601 20417 611
rect 20541 601 20575 611
rect 20263 600 20365 601
rect 20383 600 20575 601
rect 20291 572 20337 573
rect 20383 319 20417 600
rect 20427 573 20451 577
rect 20507 573 20531 577
rect 20421 572 20467 573
rect 20427 353 20451 572
rect 20459 369 20461 561
rect 20463 400 20467 572
rect 20485 572 20537 573
rect 20485 357 20531 572
rect 20507 353 20531 357
rect 20541 353 20575 600
rect 20525 319 20575 353
rect 20343 285 20359 319
rect 20383 269 20415 319
rect 20543 269 20575 319
rect 20383 258 20394 269
rect 20549 217 20575 269
rect 20583 661 20617 713
rect 20749 679 20775 713
rect 20583 611 20615 661
rect 20725 651 20775 679
rect 20725 645 20741 651
rect 20743 611 20775 651
rect 20583 601 20617 611
rect 20741 601 20775 611
rect 20583 600 20775 601
rect 20583 319 20617 600
rect 20627 573 20651 577
rect 20707 573 20731 577
rect 20621 572 20667 573
rect 20627 353 20651 572
rect 20659 369 20661 561
rect 20663 400 20667 572
rect 20685 572 20737 573
rect 20685 357 20731 572
rect 20707 353 20731 357
rect 20741 353 20775 600
rect 20725 319 20775 353
rect 20583 269 20615 319
rect 20743 269 20775 319
rect 20583 217 20617 269
rect 20749 217 20775 269
rect 20783 661 20817 713
rect 20949 679 20975 713
rect 20783 611 20815 661
rect 20925 651 20975 679
rect 20925 645 20941 651
rect 20943 611 20975 651
rect 20783 601 20817 611
rect 20941 601 20975 611
rect 20783 600 20975 601
rect 20783 319 20817 600
rect 20827 573 20851 577
rect 20907 573 20931 577
rect 20821 572 20867 573
rect 20827 353 20851 572
rect 20859 369 20861 561
rect 20863 400 20867 572
rect 20885 572 20937 573
rect 20885 357 20931 572
rect 20907 353 20931 357
rect 20941 353 20975 600
rect 20925 319 20975 353
rect 20783 269 20815 319
rect 20943 269 20975 319
rect 20783 217 20817 269
rect 20949 217 20975 269
rect 20983 661 21017 713
rect 21149 679 21175 713
rect 20983 611 21015 661
rect 21125 651 21175 679
rect 21125 645 21141 651
rect 21143 611 21175 651
rect 20983 601 21017 611
rect 21141 601 21175 611
rect 20983 600 21175 601
rect 20983 319 21017 600
rect 21027 573 21051 577
rect 21107 573 21131 577
rect 21021 572 21067 573
rect 21027 353 21051 572
rect 21059 369 21061 561
rect 21063 400 21067 572
rect 21085 572 21137 573
rect 21085 357 21131 572
rect 21107 353 21131 357
rect 21141 353 21175 600
rect 21125 319 21175 353
rect 20983 269 21015 319
rect 21143 269 21175 319
rect 20983 217 21017 269
rect 21149 217 21175 269
rect 21183 661 21217 713
rect 21183 611 21215 661
rect 21325 651 21375 679
rect 21325 645 21341 651
rect 21343 611 21375 651
rect 21399 611 21409 645
rect 21183 601 21217 611
rect 21341 601 21375 611
rect 21183 600 21375 601
rect 21393 600 21495 601
rect 21183 319 21217 600
rect 21227 573 21251 577
rect 21307 573 21331 577
rect 21221 572 21267 573
rect 21227 353 21251 572
rect 21259 369 21261 561
rect 21263 400 21267 572
rect 21285 572 21337 573
rect 21285 357 21331 572
rect 21307 353 21331 357
rect 21341 353 21375 600
rect 21421 572 21467 573
rect 21325 319 21375 353
rect 21183 269 21215 319
rect 21343 269 21375 319
rect 21399 285 21409 319
rect 21183 217 21217 269
rect 21364 258 21375 269
rect 21547 217 21617 731
rect 21947 713 22029 747
rect 22079 713 23279 747
rect 23347 731 23429 749
rect 23729 747 23812 749
rect 25147 765 25211 783
rect 25547 765 25612 783
rect 25147 749 25612 765
rect 21663 600 21765 610
rect 21793 600 21895 610
rect 21691 572 21737 582
rect 21821 572 21867 582
rect 21947 217 22017 713
rect 22349 679 22375 713
rect 22183 661 22194 672
rect 22143 611 22159 645
rect 22183 611 22215 661
rect 22325 651 22375 679
rect 22325 645 22341 651
rect 22343 611 22375 651
rect 22183 601 22217 611
rect 22341 601 22375 611
rect 22063 600 22165 601
rect 22183 600 22375 601
rect 22091 572 22137 573
rect 22183 319 22217 600
rect 22227 573 22251 577
rect 22307 573 22331 577
rect 22221 572 22267 573
rect 22227 353 22251 572
rect 22259 369 22261 561
rect 22263 400 22267 572
rect 22285 572 22337 573
rect 22285 357 22331 572
rect 22307 353 22331 357
rect 22341 353 22375 600
rect 22325 319 22375 353
rect 22143 285 22159 319
rect 22183 269 22215 319
rect 22343 269 22375 319
rect 22183 258 22194 269
rect 22349 217 22375 269
rect 22383 661 22417 713
rect 22549 679 22575 713
rect 22383 611 22415 661
rect 22525 651 22575 679
rect 22525 645 22541 651
rect 22543 611 22575 651
rect 22383 601 22417 611
rect 22541 601 22575 611
rect 22383 600 22575 601
rect 22383 319 22417 600
rect 22427 573 22451 577
rect 22507 573 22531 577
rect 22421 572 22467 573
rect 22427 353 22451 572
rect 22459 369 22461 561
rect 22463 400 22467 572
rect 22485 572 22537 573
rect 22485 357 22531 572
rect 22507 353 22531 357
rect 22541 353 22575 600
rect 22525 319 22575 353
rect 22383 269 22415 319
rect 22543 269 22575 319
rect 22383 217 22417 269
rect 22549 217 22575 269
rect 22583 661 22617 713
rect 22749 679 22775 713
rect 22583 611 22615 661
rect 22725 651 22775 679
rect 22725 645 22741 651
rect 22743 611 22775 651
rect 22583 601 22617 611
rect 22741 601 22775 611
rect 22583 600 22775 601
rect 22583 319 22617 600
rect 22627 573 22651 577
rect 22707 573 22731 577
rect 22621 572 22667 573
rect 22627 353 22651 572
rect 22659 369 22661 561
rect 22663 400 22667 572
rect 22685 572 22737 573
rect 22685 357 22731 572
rect 22707 353 22731 357
rect 22741 353 22775 600
rect 22725 319 22775 353
rect 22583 269 22615 319
rect 22743 269 22775 319
rect 22583 217 22617 269
rect 22749 217 22775 269
rect 22783 661 22817 713
rect 22949 679 22975 713
rect 22783 611 22815 661
rect 22925 651 22975 679
rect 22925 645 22941 651
rect 22943 611 22975 651
rect 22783 601 22817 611
rect 22941 601 22975 611
rect 22783 600 22975 601
rect 22783 319 22817 600
rect 22827 573 22851 577
rect 22907 573 22931 577
rect 22821 572 22867 573
rect 22827 353 22851 572
rect 22859 369 22861 561
rect 22863 400 22867 572
rect 22885 572 22937 573
rect 22885 357 22931 572
rect 22907 353 22931 357
rect 22941 353 22975 600
rect 22925 319 22975 353
rect 22783 269 22815 319
rect 22943 269 22975 319
rect 22783 217 22817 269
rect 22949 217 22975 269
rect 22983 661 23017 713
rect 22983 611 23015 661
rect 23125 651 23175 679
rect 23125 645 23141 651
rect 23143 611 23175 651
rect 23199 611 23209 645
rect 22983 601 23017 611
rect 23141 601 23175 611
rect 22983 600 23175 601
rect 23193 600 23295 601
rect 22983 319 23017 600
rect 23027 573 23051 577
rect 23107 573 23131 577
rect 23021 572 23067 573
rect 23027 353 23051 572
rect 23059 369 23061 561
rect 23063 400 23067 572
rect 23085 572 23137 573
rect 23085 357 23131 572
rect 23107 353 23131 357
rect 23141 353 23175 600
rect 23221 572 23267 573
rect 23125 319 23175 353
rect 22983 269 23015 319
rect 23143 269 23175 319
rect 23199 285 23209 319
rect 22983 217 23017 269
rect 23164 258 23175 269
rect 23347 217 23417 731
rect 23747 713 23829 747
rect 23879 713 25079 747
rect 25147 731 25229 749
rect 25529 747 25612 749
rect 26947 765 27011 783
rect 27347 765 27412 783
rect 26947 749 27412 765
rect 23463 600 23565 610
rect 23593 600 23695 610
rect 23491 572 23537 582
rect 23621 572 23667 582
rect 23747 217 23817 713
rect 24149 679 24175 713
rect 23983 661 23994 672
rect 23943 611 23959 645
rect 23983 611 24015 661
rect 24125 651 24175 679
rect 24125 645 24141 651
rect 24143 611 24175 651
rect 23983 601 24017 611
rect 24141 601 24175 611
rect 23863 600 23965 601
rect 23983 600 24175 601
rect 23891 572 23937 573
rect 23983 319 24017 600
rect 24027 573 24051 577
rect 24107 573 24131 577
rect 24021 572 24067 573
rect 24027 353 24051 572
rect 24059 369 24061 561
rect 24063 400 24067 572
rect 24085 572 24137 573
rect 24085 357 24131 572
rect 24107 353 24131 357
rect 24141 353 24175 600
rect 24125 319 24175 353
rect 23943 285 23959 319
rect 23983 269 24015 319
rect 24143 269 24175 319
rect 23983 258 23994 269
rect 24149 217 24175 269
rect 24183 661 24217 713
rect 24349 679 24375 713
rect 24183 611 24215 661
rect 24325 651 24375 679
rect 24325 645 24341 651
rect 24343 611 24375 651
rect 24183 601 24217 611
rect 24341 601 24375 611
rect 24183 600 24375 601
rect 24183 319 24217 600
rect 24227 573 24251 577
rect 24307 573 24331 577
rect 24221 572 24267 573
rect 24227 353 24251 572
rect 24259 369 24261 561
rect 24263 400 24267 572
rect 24285 572 24337 573
rect 24285 357 24331 572
rect 24307 353 24331 357
rect 24341 353 24375 600
rect 24325 319 24375 353
rect 24183 269 24215 319
rect 24343 269 24375 319
rect 24183 217 24217 269
rect 24349 217 24375 269
rect 24383 661 24417 713
rect 24549 679 24575 713
rect 24383 611 24415 661
rect 24525 651 24575 679
rect 24525 645 24541 651
rect 24543 611 24575 651
rect 24383 601 24417 611
rect 24541 601 24575 611
rect 24383 600 24575 601
rect 24383 319 24417 600
rect 24427 573 24451 577
rect 24507 573 24531 577
rect 24421 572 24467 573
rect 24427 353 24451 572
rect 24459 369 24461 561
rect 24463 400 24467 572
rect 24485 572 24537 573
rect 24485 357 24531 572
rect 24507 353 24531 357
rect 24541 353 24575 600
rect 24525 319 24575 353
rect 24383 269 24415 319
rect 24543 269 24575 319
rect 24383 217 24417 269
rect 24549 217 24575 269
rect 24583 661 24617 713
rect 24749 679 24775 713
rect 24583 611 24615 661
rect 24725 651 24775 679
rect 24725 645 24741 651
rect 24743 611 24775 651
rect 24583 601 24617 611
rect 24741 601 24775 611
rect 24583 600 24775 601
rect 24583 319 24617 600
rect 24627 573 24651 577
rect 24707 573 24731 577
rect 24621 572 24667 573
rect 24627 353 24651 572
rect 24659 369 24661 561
rect 24663 400 24667 572
rect 24685 572 24737 573
rect 24685 357 24731 572
rect 24707 353 24731 357
rect 24741 353 24775 600
rect 24725 319 24775 353
rect 24583 269 24615 319
rect 24743 269 24775 319
rect 24583 217 24617 269
rect 24749 217 24775 269
rect 24783 661 24817 713
rect 24783 611 24815 661
rect 24925 651 24975 679
rect 24925 645 24941 651
rect 24943 611 24975 651
rect 24999 611 25009 645
rect 24783 601 24817 611
rect 24941 601 24975 611
rect 24783 600 24975 601
rect 24993 600 25095 601
rect 24783 319 24817 600
rect 24827 573 24851 577
rect 24907 573 24931 577
rect 24821 572 24867 573
rect 24827 353 24851 572
rect 24859 369 24861 561
rect 24863 400 24867 572
rect 24885 572 24937 573
rect 24885 357 24931 572
rect 24907 353 24931 357
rect 24941 353 24975 600
rect 25021 572 25067 573
rect 24925 319 24975 353
rect 24783 269 24815 319
rect 24943 269 24975 319
rect 24999 285 25009 319
rect 24783 217 24817 269
rect 24964 258 24975 269
rect 25147 217 25217 731
rect 25547 713 25629 747
rect 25679 713 26879 747
rect 26947 731 27029 749
rect 27329 747 27412 749
rect 28747 765 28811 783
rect 29147 765 29212 783
rect 28747 749 29212 765
rect 25263 600 25365 610
rect 25393 600 25495 610
rect 25291 572 25337 582
rect 25421 572 25467 582
rect 25547 217 25617 713
rect 25949 679 25975 713
rect 25783 661 25794 672
rect 25743 611 25759 645
rect 25783 611 25815 661
rect 25925 651 25975 679
rect 25925 645 25941 651
rect 25943 611 25975 651
rect 25783 601 25817 611
rect 25941 601 25975 611
rect 25663 600 25765 601
rect 25783 600 25975 601
rect 25691 572 25737 573
rect 25783 319 25817 600
rect 25827 573 25851 577
rect 25907 573 25931 577
rect 25821 572 25867 573
rect 25827 353 25851 572
rect 25859 369 25861 561
rect 25863 400 25867 572
rect 25885 572 25937 573
rect 25885 357 25931 572
rect 25907 353 25931 357
rect 25941 353 25975 600
rect 25925 319 25975 353
rect 25743 285 25759 319
rect 25783 269 25815 319
rect 25943 269 25975 319
rect 25783 258 25794 269
rect 25949 217 25975 269
rect 25983 661 26017 713
rect 26149 679 26175 713
rect 25983 611 26015 661
rect 26125 651 26175 679
rect 26125 645 26141 651
rect 26143 611 26175 651
rect 25983 601 26017 611
rect 26141 601 26175 611
rect 25983 600 26175 601
rect 25983 319 26017 600
rect 26027 573 26051 577
rect 26107 573 26131 577
rect 26021 572 26067 573
rect 26027 353 26051 572
rect 26059 369 26061 561
rect 26063 400 26067 572
rect 26085 572 26137 573
rect 26085 357 26131 572
rect 26107 353 26131 357
rect 26141 353 26175 600
rect 26125 319 26175 353
rect 25983 269 26015 319
rect 26143 269 26175 319
rect 25983 217 26017 269
rect 26149 217 26175 269
rect 26183 661 26217 713
rect 26349 679 26375 713
rect 26183 611 26215 661
rect 26325 651 26375 679
rect 26325 645 26341 651
rect 26343 611 26375 651
rect 26183 601 26217 611
rect 26341 601 26375 611
rect 26183 600 26375 601
rect 26183 319 26217 600
rect 26227 573 26251 577
rect 26307 573 26331 577
rect 26221 572 26267 573
rect 26227 353 26251 572
rect 26259 369 26261 561
rect 26263 400 26267 572
rect 26285 572 26337 573
rect 26285 357 26331 572
rect 26307 353 26331 357
rect 26341 353 26375 600
rect 26325 319 26375 353
rect 26183 269 26215 319
rect 26343 269 26375 319
rect 26183 217 26217 269
rect 26349 217 26375 269
rect 26383 661 26417 713
rect 26549 679 26575 713
rect 26383 611 26415 661
rect 26525 651 26575 679
rect 26525 645 26541 651
rect 26543 611 26575 651
rect 26383 601 26417 611
rect 26541 601 26575 611
rect 26383 600 26575 601
rect 26383 319 26417 600
rect 26427 573 26451 577
rect 26507 573 26531 577
rect 26421 572 26467 573
rect 26427 353 26451 572
rect 26459 369 26461 561
rect 26463 400 26467 572
rect 26485 572 26537 573
rect 26485 357 26531 572
rect 26507 353 26531 357
rect 26541 353 26575 600
rect 26525 319 26575 353
rect 26383 269 26415 319
rect 26543 269 26575 319
rect 26383 217 26417 269
rect 26549 217 26575 269
rect 26583 661 26617 713
rect 26583 611 26615 661
rect 26725 651 26775 679
rect 26725 645 26741 651
rect 26743 611 26775 651
rect 26799 611 26809 645
rect 26583 601 26617 611
rect 26741 601 26775 611
rect 26583 600 26775 601
rect 26793 600 26895 601
rect 26583 319 26617 600
rect 26627 573 26651 577
rect 26707 573 26731 577
rect 26621 572 26667 573
rect 26627 353 26651 572
rect 26659 369 26661 561
rect 26663 400 26667 572
rect 26685 572 26737 573
rect 26685 357 26731 572
rect 26707 353 26731 357
rect 26741 353 26775 600
rect 26821 572 26867 573
rect 26725 319 26775 353
rect 26583 269 26615 319
rect 26743 269 26775 319
rect 26799 285 26809 319
rect 26583 217 26617 269
rect 26764 258 26775 269
rect 26947 217 27017 731
rect 27347 713 27429 747
rect 27479 713 28679 747
rect 28747 731 28829 749
rect 29129 747 29212 749
rect 30547 765 30611 783
rect 30947 765 31012 783
rect 30547 749 31012 765
rect 27063 600 27165 610
rect 27193 600 27295 610
rect 27091 572 27137 582
rect 27221 572 27267 582
rect 27347 217 27417 713
rect 27749 679 27775 713
rect 27583 661 27594 672
rect 27543 611 27559 645
rect 27583 611 27615 661
rect 27725 651 27775 679
rect 27725 645 27741 651
rect 27743 611 27775 651
rect 27583 601 27617 611
rect 27741 601 27775 611
rect 27463 600 27565 601
rect 27583 600 27775 601
rect 27491 572 27537 573
rect 27583 319 27617 600
rect 27627 573 27651 577
rect 27707 573 27731 577
rect 27621 572 27667 573
rect 27627 353 27651 572
rect 27659 369 27661 561
rect 27663 400 27667 572
rect 27685 572 27737 573
rect 27685 357 27731 572
rect 27707 353 27731 357
rect 27741 353 27775 600
rect 27725 319 27775 353
rect 27543 285 27559 319
rect 27583 269 27615 319
rect 27743 269 27775 319
rect 27583 258 27594 269
rect 27749 217 27775 269
rect 27783 661 27817 713
rect 27949 679 27975 713
rect 27783 611 27815 661
rect 27925 651 27975 679
rect 27925 645 27941 651
rect 27943 611 27975 651
rect 27783 601 27817 611
rect 27941 601 27975 611
rect 27783 600 27975 601
rect 27783 319 27817 600
rect 27827 573 27851 577
rect 27907 573 27931 577
rect 27821 572 27867 573
rect 27827 353 27851 572
rect 27859 369 27861 561
rect 27863 400 27867 572
rect 27885 572 27937 573
rect 27885 357 27931 572
rect 27907 353 27931 357
rect 27941 353 27975 600
rect 27925 319 27975 353
rect 27783 269 27815 319
rect 27943 269 27975 319
rect 27783 217 27817 269
rect 27949 217 27975 269
rect 27983 661 28017 713
rect 28149 679 28175 713
rect 27983 611 28015 661
rect 28125 651 28175 679
rect 28125 645 28141 651
rect 28143 611 28175 651
rect 27983 601 28017 611
rect 28141 601 28175 611
rect 27983 600 28175 601
rect 27983 319 28017 600
rect 28027 573 28051 577
rect 28107 573 28131 577
rect 28021 572 28067 573
rect 28027 353 28051 572
rect 28059 369 28061 561
rect 28063 400 28067 572
rect 28085 572 28137 573
rect 28085 357 28131 572
rect 28107 353 28131 357
rect 28141 353 28175 600
rect 28125 319 28175 353
rect 27983 269 28015 319
rect 28143 269 28175 319
rect 27983 217 28017 269
rect 28149 217 28175 269
rect 28183 661 28217 713
rect 28349 679 28375 713
rect 28183 611 28215 661
rect 28325 651 28375 679
rect 28325 645 28341 651
rect 28343 611 28375 651
rect 28183 601 28217 611
rect 28341 601 28375 611
rect 28183 600 28375 601
rect 28183 319 28217 600
rect 28227 573 28251 577
rect 28307 573 28331 577
rect 28221 572 28267 573
rect 28227 353 28251 572
rect 28259 369 28261 561
rect 28263 400 28267 572
rect 28285 572 28337 573
rect 28285 357 28331 572
rect 28307 353 28331 357
rect 28341 353 28375 600
rect 28325 319 28375 353
rect 28183 269 28215 319
rect 28343 269 28375 319
rect 28183 217 28217 269
rect 28349 217 28375 269
rect 28383 661 28417 713
rect 28383 611 28415 661
rect 28525 651 28575 679
rect 28525 645 28541 651
rect 28543 611 28575 651
rect 28599 611 28609 645
rect 28383 601 28417 611
rect 28541 601 28575 611
rect 28383 600 28575 601
rect 28593 600 28695 601
rect 28383 319 28417 600
rect 28427 573 28451 577
rect 28507 573 28531 577
rect 28421 572 28467 573
rect 28427 353 28451 572
rect 28459 369 28461 561
rect 28463 400 28467 572
rect 28485 572 28537 573
rect 28485 357 28531 572
rect 28507 353 28531 357
rect 28541 353 28575 600
rect 28621 572 28667 573
rect 28525 319 28575 353
rect 28383 269 28415 319
rect 28543 269 28575 319
rect 28599 285 28609 319
rect 28383 217 28417 269
rect 28564 258 28575 269
rect 28747 217 28817 731
rect 29147 713 29229 747
rect 29279 713 30479 747
rect 30547 731 30629 749
rect 30929 747 31012 749
rect 32347 765 32411 783
rect 32747 765 32812 783
rect 32347 749 32812 765
rect 28863 600 28965 610
rect 28993 600 29095 610
rect 28891 572 28937 582
rect 29021 572 29067 582
rect 29147 217 29217 713
rect 29549 679 29575 713
rect 29383 661 29394 672
rect 29343 611 29359 645
rect 29383 611 29415 661
rect 29525 651 29575 679
rect 29525 645 29541 651
rect 29543 611 29575 651
rect 29383 601 29417 611
rect 29541 601 29575 611
rect 29263 600 29365 601
rect 29383 600 29575 601
rect 29291 572 29337 573
rect 29383 319 29417 600
rect 29427 573 29451 577
rect 29507 573 29531 577
rect 29421 572 29467 573
rect 29427 353 29451 572
rect 29459 369 29461 561
rect 29463 400 29467 572
rect 29485 572 29537 573
rect 29485 357 29531 572
rect 29507 353 29531 357
rect 29541 353 29575 600
rect 29525 319 29575 353
rect 29343 285 29359 319
rect 29383 269 29415 319
rect 29543 269 29575 319
rect 29383 258 29394 269
rect 29549 217 29575 269
rect 29583 661 29617 713
rect 29749 679 29775 713
rect 29583 611 29615 661
rect 29725 651 29775 679
rect 29725 645 29741 651
rect 29743 611 29775 651
rect 29583 601 29617 611
rect 29741 601 29775 611
rect 29583 600 29775 601
rect 29583 319 29617 600
rect 29627 573 29651 577
rect 29707 573 29731 577
rect 29621 572 29667 573
rect 29627 353 29651 572
rect 29659 369 29661 561
rect 29663 400 29667 572
rect 29685 572 29737 573
rect 29685 357 29731 572
rect 29707 353 29731 357
rect 29741 353 29775 600
rect 29725 319 29775 353
rect 29583 269 29615 319
rect 29743 269 29775 319
rect 29583 217 29617 269
rect 29749 217 29775 269
rect 29783 661 29817 713
rect 29949 679 29975 713
rect 29783 611 29815 661
rect 29925 651 29975 679
rect 29925 645 29941 651
rect 29943 611 29975 651
rect 29783 601 29817 611
rect 29941 601 29975 611
rect 29783 600 29975 601
rect 29783 319 29817 600
rect 29827 573 29851 577
rect 29907 573 29931 577
rect 29821 572 29867 573
rect 29827 353 29851 572
rect 29859 369 29861 561
rect 29863 400 29867 572
rect 29885 572 29937 573
rect 29885 357 29931 572
rect 29907 353 29931 357
rect 29941 353 29975 600
rect 29925 319 29975 353
rect 29783 269 29815 319
rect 29943 269 29975 319
rect 29783 217 29817 269
rect 29949 217 29975 269
rect 29983 661 30017 713
rect 30149 679 30175 713
rect 29983 611 30015 661
rect 30125 651 30175 679
rect 30125 645 30141 651
rect 30143 611 30175 651
rect 29983 601 30017 611
rect 30141 601 30175 611
rect 29983 600 30175 601
rect 29983 319 30017 600
rect 30027 573 30051 577
rect 30107 573 30131 577
rect 30021 572 30067 573
rect 30027 353 30051 572
rect 30059 369 30061 561
rect 30063 400 30067 572
rect 30085 572 30137 573
rect 30085 357 30131 572
rect 30107 353 30131 357
rect 30141 353 30175 600
rect 30125 319 30175 353
rect 29983 269 30015 319
rect 30143 269 30175 319
rect 29983 217 30017 269
rect 30149 217 30175 269
rect 30183 661 30217 713
rect 30183 611 30215 661
rect 30325 651 30375 679
rect 30325 645 30341 651
rect 30343 611 30375 651
rect 30399 611 30409 645
rect 30183 601 30217 611
rect 30341 601 30375 611
rect 30183 600 30375 601
rect 30393 600 30495 601
rect 30183 319 30217 600
rect 30227 573 30251 577
rect 30307 573 30331 577
rect 30221 572 30267 573
rect 30227 353 30251 572
rect 30259 369 30261 561
rect 30263 400 30267 572
rect 30285 572 30337 573
rect 30285 357 30331 572
rect 30307 353 30331 357
rect 30341 353 30375 600
rect 30421 572 30467 573
rect 30325 319 30375 353
rect 30183 269 30215 319
rect 30343 269 30375 319
rect 30399 285 30409 319
rect 30183 217 30217 269
rect 30364 258 30375 269
rect 30547 217 30617 731
rect 30947 713 31029 747
rect 31079 713 32279 747
rect 32347 731 32429 749
rect 32729 747 32812 749
rect 34147 765 34211 783
rect 34547 765 34612 783
rect 34147 749 34612 765
rect 30663 600 30765 610
rect 30793 600 30895 610
rect 30691 572 30737 582
rect 30821 572 30867 582
rect 30947 217 31017 713
rect 31349 679 31375 713
rect 31183 661 31194 672
rect 31143 611 31159 645
rect 31183 611 31215 661
rect 31325 651 31375 679
rect 31325 645 31341 651
rect 31343 611 31375 651
rect 31183 601 31217 611
rect 31341 601 31375 611
rect 31063 600 31165 601
rect 31183 600 31375 601
rect 31091 572 31137 573
rect 31183 319 31217 600
rect 31227 573 31251 577
rect 31307 573 31331 577
rect 31221 572 31267 573
rect 31227 353 31251 572
rect 31259 369 31261 561
rect 31263 400 31267 572
rect 31285 572 31337 573
rect 31285 357 31331 572
rect 31307 353 31331 357
rect 31341 353 31375 600
rect 31325 319 31375 353
rect 31143 285 31159 319
rect 31183 269 31215 319
rect 31343 269 31375 319
rect 31183 258 31194 269
rect 31349 217 31375 269
rect 31383 661 31417 713
rect 31549 679 31575 713
rect 31383 611 31415 661
rect 31525 651 31575 679
rect 31525 645 31541 651
rect 31543 611 31575 651
rect 31383 601 31417 611
rect 31541 601 31575 611
rect 31383 600 31575 601
rect 31383 319 31417 600
rect 31427 573 31451 577
rect 31507 573 31531 577
rect 31421 572 31467 573
rect 31427 353 31451 572
rect 31459 369 31461 561
rect 31463 400 31467 572
rect 31485 572 31537 573
rect 31485 357 31531 572
rect 31507 353 31531 357
rect 31541 353 31575 600
rect 31525 319 31575 353
rect 31383 269 31415 319
rect 31543 269 31575 319
rect 31383 217 31417 269
rect 31549 217 31575 269
rect 31583 661 31617 713
rect 31749 679 31775 713
rect 31583 611 31615 661
rect 31725 651 31775 679
rect 31725 645 31741 651
rect 31743 611 31775 651
rect 31583 601 31617 611
rect 31741 601 31775 611
rect 31583 600 31775 601
rect 31583 319 31617 600
rect 31627 573 31651 577
rect 31707 573 31731 577
rect 31621 572 31667 573
rect 31627 353 31651 572
rect 31659 369 31661 561
rect 31663 400 31667 572
rect 31685 572 31737 573
rect 31685 357 31731 572
rect 31707 353 31731 357
rect 31741 353 31775 600
rect 31725 319 31775 353
rect 31583 269 31615 319
rect 31743 269 31775 319
rect 31583 217 31617 269
rect 31749 217 31775 269
rect 31783 661 31817 713
rect 31949 679 31975 713
rect 31783 611 31815 661
rect 31925 651 31975 679
rect 31925 645 31941 651
rect 31943 611 31975 651
rect 31783 601 31817 611
rect 31941 601 31975 611
rect 31783 600 31975 601
rect 31783 319 31817 600
rect 31827 573 31851 577
rect 31907 573 31931 577
rect 31821 572 31867 573
rect 31827 353 31851 572
rect 31859 369 31861 561
rect 31863 400 31867 572
rect 31885 572 31937 573
rect 31885 357 31931 572
rect 31907 353 31931 357
rect 31941 353 31975 600
rect 31925 319 31975 353
rect 31783 269 31815 319
rect 31943 269 31975 319
rect 31783 217 31817 269
rect 31949 217 31975 269
rect 31983 661 32017 713
rect 31983 611 32015 661
rect 32125 651 32175 679
rect 32125 645 32141 651
rect 32143 611 32175 651
rect 32199 611 32209 645
rect 31983 601 32017 611
rect 32141 601 32175 611
rect 31983 600 32175 601
rect 32193 600 32295 601
rect 31983 319 32017 600
rect 32027 573 32051 577
rect 32107 573 32131 577
rect 32021 572 32067 573
rect 32027 353 32051 572
rect 32059 369 32061 561
rect 32063 400 32067 572
rect 32085 572 32137 573
rect 32085 357 32131 572
rect 32107 353 32131 357
rect 32141 353 32175 600
rect 32221 572 32267 573
rect 32125 319 32175 353
rect 31983 269 32015 319
rect 32143 269 32175 319
rect 32199 285 32209 319
rect 31983 217 32017 269
rect 32164 258 32175 269
rect 32347 217 32417 731
rect 32747 713 32829 747
rect 32879 713 34079 747
rect 34147 731 34229 749
rect 34529 747 34612 749
rect 35947 765 36011 783
rect 36347 765 36412 783
rect 35947 749 36412 765
rect 32463 600 32565 610
rect 32593 600 32695 610
rect 32491 572 32537 582
rect 32621 572 32667 582
rect 32747 217 32817 713
rect 33149 679 33175 713
rect 32983 661 32994 672
rect 32943 611 32959 645
rect 32983 611 33015 661
rect 33125 651 33175 679
rect 33125 645 33141 651
rect 33143 611 33175 651
rect 32983 601 33017 611
rect 33141 601 33175 611
rect 32863 600 32965 601
rect 32983 600 33175 601
rect 32891 572 32937 573
rect 32983 319 33017 600
rect 33027 573 33051 577
rect 33107 573 33131 577
rect 33021 572 33067 573
rect 33027 353 33051 572
rect 33059 369 33061 561
rect 33063 400 33067 572
rect 33085 572 33137 573
rect 33085 357 33131 572
rect 33107 353 33131 357
rect 33141 353 33175 600
rect 33125 319 33175 353
rect 32943 285 32959 319
rect 32983 269 33015 319
rect 33143 269 33175 319
rect 32983 258 32994 269
rect 33149 217 33175 269
rect 33183 661 33217 713
rect 33349 679 33375 713
rect 33183 611 33215 661
rect 33325 651 33375 679
rect 33325 645 33341 651
rect 33343 611 33375 651
rect 33183 601 33217 611
rect 33341 601 33375 611
rect 33183 600 33375 601
rect 33183 319 33217 600
rect 33227 573 33251 577
rect 33307 573 33331 577
rect 33221 572 33267 573
rect 33227 353 33251 572
rect 33259 369 33261 561
rect 33263 400 33267 572
rect 33285 572 33337 573
rect 33285 357 33331 572
rect 33307 353 33331 357
rect 33341 353 33375 600
rect 33325 319 33375 353
rect 33183 269 33215 319
rect 33343 269 33375 319
rect 33183 217 33217 269
rect 33349 217 33375 269
rect 33383 661 33417 713
rect 33549 679 33575 713
rect 33383 611 33415 661
rect 33525 651 33575 679
rect 33525 645 33541 651
rect 33543 611 33575 651
rect 33383 601 33417 611
rect 33541 601 33575 611
rect 33383 600 33575 601
rect 33383 319 33417 600
rect 33427 573 33451 577
rect 33507 573 33531 577
rect 33421 572 33467 573
rect 33427 353 33451 572
rect 33459 369 33461 561
rect 33463 400 33467 572
rect 33485 572 33537 573
rect 33485 357 33531 572
rect 33507 353 33531 357
rect 33541 353 33575 600
rect 33525 319 33575 353
rect 33383 269 33415 319
rect 33543 269 33575 319
rect 33383 217 33417 269
rect 33549 217 33575 269
rect 33583 661 33617 713
rect 33749 679 33775 713
rect 33583 611 33615 661
rect 33725 651 33775 679
rect 33725 645 33741 651
rect 33743 611 33775 651
rect 33583 601 33617 611
rect 33741 601 33775 611
rect 33583 600 33775 601
rect 33583 319 33617 600
rect 33627 573 33651 577
rect 33707 573 33731 577
rect 33621 572 33667 573
rect 33627 353 33651 572
rect 33659 369 33661 561
rect 33663 400 33667 572
rect 33685 572 33737 573
rect 33685 357 33731 572
rect 33707 353 33731 357
rect 33741 353 33775 600
rect 33725 319 33775 353
rect 33583 269 33615 319
rect 33743 269 33775 319
rect 33583 217 33617 269
rect 33749 217 33775 269
rect 33783 661 33817 713
rect 33783 611 33815 661
rect 33925 651 33975 679
rect 33925 645 33941 651
rect 33943 611 33975 651
rect 33999 611 34009 645
rect 33783 601 33817 611
rect 33941 601 33975 611
rect 33783 600 33975 601
rect 33993 600 34095 601
rect 33783 319 33817 600
rect 33827 573 33851 577
rect 33907 573 33931 577
rect 33821 572 33867 573
rect 33827 353 33851 572
rect 33859 369 33861 561
rect 33863 400 33867 572
rect 33885 572 33937 573
rect 33885 357 33931 572
rect 33907 353 33931 357
rect 33941 353 33975 600
rect 34021 572 34067 573
rect 33925 319 33975 353
rect 33783 269 33815 319
rect 33943 269 33975 319
rect 33999 285 34009 319
rect 33783 217 33817 269
rect 33964 258 33975 269
rect 34147 217 34217 731
rect 34547 713 34629 747
rect 34679 713 35879 747
rect 35947 731 36029 749
rect 36329 747 36412 749
rect 37747 765 37811 783
rect 38147 765 38212 783
rect 37747 749 38212 765
rect 34263 600 34365 610
rect 34393 600 34495 610
rect 34291 572 34337 582
rect 34421 572 34467 582
rect 34547 217 34617 713
rect 34949 679 34975 713
rect 34783 661 34794 672
rect 34743 611 34759 645
rect 34783 611 34815 661
rect 34925 651 34975 679
rect 34925 645 34941 651
rect 34943 611 34975 651
rect 34783 601 34817 611
rect 34941 601 34975 611
rect 34663 600 34765 601
rect 34783 600 34975 601
rect 34691 572 34737 573
rect 34783 319 34817 600
rect 34827 573 34851 577
rect 34907 573 34931 577
rect 34821 572 34867 573
rect 34827 353 34851 572
rect 34859 369 34861 561
rect 34863 400 34867 572
rect 34885 572 34937 573
rect 34885 357 34931 572
rect 34907 353 34931 357
rect 34941 353 34975 600
rect 34925 319 34975 353
rect 34743 285 34759 319
rect 34783 269 34815 319
rect 34943 269 34975 319
rect 34783 258 34794 269
rect 34949 217 34975 269
rect 34983 661 35017 713
rect 35149 679 35175 713
rect 34983 611 35015 661
rect 35125 651 35175 679
rect 35125 645 35141 651
rect 35143 611 35175 651
rect 34983 601 35017 611
rect 35141 601 35175 611
rect 34983 600 35175 601
rect 34983 319 35017 600
rect 35027 573 35051 577
rect 35107 573 35131 577
rect 35021 572 35067 573
rect 35027 353 35051 572
rect 35059 369 35061 561
rect 35063 400 35067 572
rect 35085 572 35137 573
rect 35085 357 35131 572
rect 35107 353 35131 357
rect 35141 353 35175 600
rect 35125 319 35175 353
rect 34983 269 35015 319
rect 35143 269 35175 319
rect 34983 217 35017 269
rect 35149 217 35175 269
rect 35183 661 35217 713
rect 35349 679 35375 713
rect 35183 611 35215 661
rect 35325 651 35375 679
rect 35325 645 35341 651
rect 35343 611 35375 651
rect 35183 601 35217 611
rect 35341 601 35375 611
rect 35183 600 35375 601
rect 35183 319 35217 600
rect 35227 573 35251 577
rect 35307 573 35331 577
rect 35221 572 35267 573
rect 35227 353 35251 572
rect 35259 369 35261 561
rect 35263 400 35267 572
rect 35285 572 35337 573
rect 35285 357 35331 572
rect 35307 353 35331 357
rect 35341 353 35375 600
rect 35325 319 35375 353
rect 35183 269 35215 319
rect 35343 269 35375 319
rect 35183 217 35217 269
rect 35349 217 35375 269
rect 35383 661 35417 713
rect 35549 679 35575 713
rect 35383 611 35415 661
rect 35525 651 35575 679
rect 35525 645 35541 651
rect 35543 611 35575 651
rect 35383 601 35417 611
rect 35541 601 35575 611
rect 35383 600 35575 601
rect 35383 319 35417 600
rect 35427 573 35451 577
rect 35507 573 35531 577
rect 35421 572 35467 573
rect 35427 353 35451 572
rect 35459 369 35461 561
rect 35463 400 35467 572
rect 35485 572 35537 573
rect 35485 357 35531 572
rect 35507 353 35531 357
rect 35541 353 35575 600
rect 35525 319 35575 353
rect 35383 269 35415 319
rect 35543 269 35575 319
rect 35383 217 35417 269
rect 35549 217 35575 269
rect 35583 661 35617 713
rect 35583 611 35615 661
rect 35725 651 35775 679
rect 35725 645 35741 651
rect 35743 611 35775 651
rect 35799 611 35809 645
rect 35583 601 35617 611
rect 35741 601 35775 611
rect 35583 600 35775 601
rect 35793 600 35895 601
rect 35583 319 35617 600
rect 35627 573 35651 577
rect 35707 573 35731 577
rect 35621 572 35667 573
rect 35627 353 35651 572
rect 35659 369 35661 561
rect 35663 400 35667 572
rect 35685 572 35737 573
rect 35685 357 35731 572
rect 35707 353 35731 357
rect 35741 353 35775 600
rect 35821 572 35867 573
rect 35725 319 35775 353
rect 35583 269 35615 319
rect 35743 269 35775 319
rect 35799 285 35809 319
rect 35583 217 35617 269
rect 35764 258 35775 269
rect 35947 217 36017 731
rect 36347 713 36429 747
rect 36479 713 37679 747
rect 37747 731 37829 749
rect 38129 747 38212 749
rect 39547 765 39611 783
rect 39947 765 40012 783
rect 39547 749 40012 765
rect 36063 600 36165 610
rect 36193 600 36295 610
rect 36091 572 36137 582
rect 36221 572 36267 582
rect 36347 217 36417 713
rect 36749 679 36775 713
rect 36583 661 36594 672
rect 36543 611 36559 645
rect 36583 611 36615 661
rect 36725 651 36775 679
rect 36725 645 36741 651
rect 36743 611 36775 651
rect 36583 601 36617 611
rect 36741 601 36775 611
rect 36463 600 36565 601
rect 36583 600 36775 601
rect 36491 572 36537 573
rect 36583 319 36617 600
rect 36627 573 36651 577
rect 36707 573 36731 577
rect 36621 572 36667 573
rect 36627 353 36651 572
rect 36659 369 36661 561
rect 36663 400 36667 572
rect 36685 572 36737 573
rect 36685 357 36731 572
rect 36707 353 36731 357
rect 36741 353 36775 600
rect 36725 319 36775 353
rect 36543 285 36559 319
rect 36583 269 36615 319
rect 36743 269 36775 319
rect 36583 258 36594 269
rect 36749 217 36775 269
rect 36783 661 36817 713
rect 36949 679 36975 713
rect 36783 611 36815 661
rect 36925 651 36975 679
rect 36925 645 36941 651
rect 36943 611 36975 651
rect 36783 601 36817 611
rect 36941 601 36975 611
rect 36783 600 36975 601
rect 36783 319 36817 600
rect 36827 573 36851 577
rect 36907 573 36931 577
rect 36821 572 36867 573
rect 36827 353 36851 572
rect 36859 369 36861 561
rect 36863 400 36867 572
rect 36885 572 36937 573
rect 36885 357 36931 572
rect 36907 353 36931 357
rect 36941 353 36975 600
rect 36925 319 36975 353
rect 36783 269 36815 319
rect 36943 269 36975 319
rect 36783 217 36817 269
rect 36949 217 36975 269
rect 36983 661 37017 713
rect 37149 679 37175 713
rect 36983 611 37015 661
rect 37125 651 37175 679
rect 37125 645 37141 651
rect 37143 611 37175 651
rect 36983 601 37017 611
rect 37141 601 37175 611
rect 36983 600 37175 601
rect 36983 319 37017 600
rect 37027 573 37051 577
rect 37107 573 37131 577
rect 37021 572 37067 573
rect 37027 353 37051 572
rect 37059 369 37061 561
rect 37063 400 37067 572
rect 37085 572 37137 573
rect 37085 357 37131 572
rect 37107 353 37131 357
rect 37141 353 37175 600
rect 37125 319 37175 353
rect 36983 269 37015 319
rect 37143 269 37175 319
rect 36983 217 37017 269
rect 37149 217 37175 269
rect 37183 661 37217 713
rect 37349 679 37375 713
rect 37183 611 37215 661
rect 37325 651 37375 679
rect 37325 645 37341 651
rect 37343 611 37375 651
rect 37183 601 37217 611
rect 37341 601 37375 611
rect 37183 600 37375 601
rect 37183 319 37217 600
rect 37227 573 37251 577
rect 37307 573 37331 577
rect 37221 572 37267 573
rect 37227 353 37251 572
rect 37259 369 37261 561
rect 37263 400 37267 572
rect 37285 572 37337 573
rect 37285 357 37331 572
rect 37307 353 37331 357
rect 37341 353 37375 600
rect 37325 319 37375 353
rect 37183 269 37215 319
rect 37343 269 37375 319
rect 37183 217 37217 269
rect 37349 217 37375 269
rect 37383 661 37417 713
rect 37383 611 37415 661
rect 37525 651 37575 679
rect 37525 645 37541 651
rect 37543 611 37575 651
rect 37599 611 37609 645
rect 37383 601 37417 611
rect 37541 601 37575 611
rect 37383 600 37575 601
rect 37593 600 37695 601
rect 37383 319 37417 600
rect 37427 573 37451 577
rect 37507 573 37531 577
rect 37421 572 37467 573
rect 37427 353 37451 572
rect 37459 369 37461 561
rect 37463 400 37467 572
rect 37485 572 37537 573
rect 37485 357 37531 572
rect 37507 353 37531 357
rect 37541 353 37575 600
rect 37621 572 37667 573
rect 37525 319 37575 353
rect 37383 269 37415 319
rect 37543 269 37575 319
rect 37599 285 37609 319
rect 37383 217 37417 269
rect 37564 258 37575 269
rect 37747 217 37817 731
rect 38147 713 38229 747
rect 38279 713 39479 747
rect 39547 731 39629 749
rect 39929 747 40012 749
rect 41347 765 41411 783
rect 41747 765 41812 783
rect 41347 749 41812 765
rect 37863 600 37965 610
rect 37993 600 38095 610
rect 37891 572 37937 582
rect 38021 572 38067 582
rect 38147 217 38217 713
rect 38549 679 38575 713
rect 38383 661 38394 672
rect 38343 611 38359 645
rect 38383 611 38415 661
rect 38525 651 38575 679
rect 38525 645 38541 651
rect 38543 611 38575 651
rect 38383 601 38417 611
rect 38541 601 38575 611
rect 38263 600 38365 601
rect 38383 600 38575 601
rect 38291 572 38337 573
rect 38383 319 38417 600
rect 38427 573 38451 577
rect 38507 573 38531 577
rect 38421 572 38467 573
rect 38427 353 38451 572
rect 38459 369 38461 561
rect 38463 400 38467 572
rect 38485 572 38537 573
rect 38485 357 38531 572
rect 38507 353 38531 357
rect 38541 353 38575 600
rect 38525 319 38575 353
rect 38343 285 38359 319
rect 38383 269 38415 319
rect 38543 269 38575 319
rect 38383 258 38394 269
rect 38549 217 38575 269
rect 38583 661 38617 713
rect 38749 679 38775 713
rect 38583 611 38615 661
rect 38725 651 38775 679
rect 38725 645 38741 651
rect 38743 611 38775 651
rect 38583 601 38617 611
rect 38741 601 38775 611
rect 38583 600 38775 601
rect 38583 319 38617 600
rect 38627 573 38651 577
rect 38707 573 38731 577
rect 38621 572 38667 573
rect 38627 353 38651 572
rect 38659 369 38661 561
rect 38663 400 38667 572
rect 38685 572 38737 573
rect 38685 357 38731 572
rect 38707 353 38731 357
rect 38741 353 38775 600
rect 38725 319 38775 353
rect 38583 269 38615 319
rect 38743 269 38775 319
rect 38583 217 38617 269
rect 38749 217 38775 269
rect 38783 661 38817 713
rect 38949 679 38975 713
rect 38783 611 38815 661
rect 38925 651 38975 679
rect 38925 645 38941 651
rect 38943 611 38975 651
rect 38783 601 38817 611
rect 38941 601 38975 611
rect 38783 600 38975 601
rect 38783 319 38817 600
rect 38827 573 38851 577
rect 38907 573 38931 577
rect 38821 572 38867 573
rect 38827 353 38851 572
rect 38859 369 38861 561
rect 38863 400 38867 572
rect 38885 572 38937 573
rect 38885 357 38931 572
rect 38907 353 38931 357
rect 38941 353 38975 600
rect 38925 319 38975 353
rect 38783 269 38815 319
rect 38943 269 38975 319
rect 38783 217 38817 269
rect 38949 217 38975 269
rect 38983 661 39017 713
rect 39149 679 39175 713
rect 38983 611 39015 661
rect 39125 651 39175 679
rect 39125 645 39141 651
rect 39143 611 39175 651
rect 38983 601 39017 611
rect 39141 601 39175 611
rect 38983 600 39175 601
rect 38983 319 39017 600
rect 39027 573 39051 577
rect 39107 573 39131 577
rect 39021 572 39067 573
rect 39027 353 39051 572
rect 39059 369 39061 561
rect 39063 400 39067 572
rect 39085 572 39137 573
rect 39085 357 39131 572
rect 39107 353 39131 357
rect 39141 353 39175 600
rect 39125 319 39175 353
rect 38983 269 39015 319
rect 39143 269 39175 319
rect 38983 217 39017 269
rect 39149 217 39175 269
rect 39183 661 39217 713
rect 39183 611 39215 661
rect 39325 651 39375 679
rect 39325 645 39341 651
rect 39343 611 39375 651
rect 39399 611 39409 645
rect 39183 601 39217 611
rect 39341 601 39375 611
rect 39183 600 39375 601
rect 39393 600 39495 601
rect 39183 319 39217 600
rect 39227 573 39251 577
rect 39307 573 39331 577
rect 39221 572 39267 573
rect 39227 353 39251 572
rect 39259 369 39261 561
rect 39263 400 39267 572
rect 39285 572 39337 573
rect 39285 357 39331 572
rect 39307 353 39331 357
rect 39341 353 39375 600
rect 39421 572 39467 573
rect 39325 319 39375 353
rect 39183 269 39215 319
rect 39343 269 39375 319
rect 39399 285 39409 319
rect 39183 217 39217 269
rect 39364 258 39375 269
rect 39547 217 39617 731
rect 39947 713 40029 747
rect 40079 713 41279 747
rect 41347 731 41429 749
rect 41729 747 41812 749
rect 43147 765 43211 783
rect 43547 765 43612 783
rect 43147 749 43612 765
rect 39663 600 39765 610
rect 39793 600 39895 610
rect 39691 572 39737 582
rect 39821 572 39867 582
rect 39947 217 40017 713
rect 40349 679 40375 713
rect 40183 661 40194 672
rect 40143 611 40159 645
rect 40183 611 40215 661
rect 40325 651 40375 679
rect 40325 645 40341 651
rect 40343 611 40375 651
rect 40183 601 40217 611
rect 40341 601 40375 611
rect 40063 600 40165 601
rect 40183 600 40375 601
rect 40091 572 40137 573
rect 40183 319 40217 600
rect 40227 573 40251 577
rect 40307 573 40331 577
rect 40221 572 40267 573
rect 40227 353 40251 572
rect 40259 369 40261 561
rect 40263 400 40267 572
rect 40285 572 40337 573
rect 40285 357 40331 572
rect 40307 353 40331 357
rect 40341 353 40375 600
rect 40325 319 40375 353
rect 40143 285 40159 319
rect 40183 269 40215 319
rect 40343 269 40375 319
rect 40183 258 40194 269
rect 40349 217 40375 269
rect 40383 661 40417 713
rect 40549 679 40575 713
rect 40383 611 40415 661
rect 40525 651 40575 679
rect 40525 645 40541 651
rect 40543 611 40575 651
rect 40383 601 40417 611
rect 40541 601 40575 611
rect 40383 600 40575 601
rect 40383 319 40417 600
rect 40427 573 40451 577
rect 40507 573 40531 577
rect 40421 572 40467 573
rect 40427 353 40451 572
rect 40459 369 40461 561
rect 40463 400 40467 572
rect 40485 572 40537 573
rect 40485 357 40531 572
rect 40507 353 40531 357
rect 40541 353 40575 600
rect 40525 319 40575 353
rect 40383 269 40415 319
rect 40543 269 40575 319
rect 40383 217 40417 269
rect 40549 217 40575 269
rect 40583 661 40617 713
rect 40749 679 40775 713
rect 40583 611 40615 661
rect 40725 651 40775 679
rect 40725 645 40741 651
rect 40743 611 40775 651
rect 40583 601 40617 611
rect 40741 601 40775 611
rect 40583 600 40775 601
rect 40583 319 40617 600
rect 40627 573 40651 577
rect 40707 573 40731 577
rect 40621 572 40667 573
rect 40627 353 40651 572
rect 40659 369 40661 561
rect 40663 400 40667 572
rect 40685 572 40737 573
rect 40685 357 40731 572
rect 40707 353 40731 357
rect 40741 353 40775 600
rect 40725 319 40775 353
rect 40583 269 40615 319
rect 40743 269 40775 319
rect 40583 217 40617 269
rect 40749 217 40775 269
rect 40783 661 40817 713
rect 40949 679 40975 713
rect 40783 611 40815 661
rect 40925 651 40975 679
rect 40925 645 40941 651
rect 40943 611 40975 651
rect 40783 601 40817 611
rect 40941 601 40975 611
rect 40783 600 40975 601
rect 40783 319 40817 600
rect 40827 573 40851 577
rect 40907 573 40931 577
rect 40821 572 40867 573
rect 40827 353 40851 572
rect 40859 369 40861 561
rect 40863 400 40867 572
rect 40885 572 40937 573
rect 40885 357 40931 572
rect 40907 353 40931 357
rect 40941 353 40975 600
rect 40925 319 40975 353
rect 40783 269 40815 319
rect 40943 269 40975 319
rect 40783 217 40817 269
rect 40949 217 40975 269
rect 40983 661 41017 713
rect 40983 611 41015 661
rect 41125 651 41175 679
rect 41125 645 41141 651
rect 41143 611 41175 651
rect 41199 611 41209 645
rect 40983 601 41017 611
rect 41141 601 41175 611
rect 40983 600 41175 601
rect 41193 600 41295 601
rect 40983 319 41017 600
rect 41027 573 41051 577
rect 41107 573 41131 577
rect 41021 572 41067 573
rect 41027 353 41051 572
rect 41059 369 41061 561
rect 41063 400 41067 572
rect 41085 572 41137 573
rect 41085 357 41131 572
rect 41107 353 41131 357
rect 41141 353 41175 600
rect 41221 572 41267 573
rect 41125 319 41175 353
rect 40983 269 41015 319
rect 41143 269 41175 319
rect 41199 285 41209 319
rect 40983 217 41017 269
rect 41164 258 41175 269
rect 41347 217 41417 731
rect 41747 713 41829 747
rect 41879 713 43079 747
rect 43147 731 43229 749
rect 43529 747 43612 749
rect 44947 765 45011 783
rect 45347 765 45412 783
rect 44947 749 45412 765
rect 41463 600 41565 610
rect 41593 600 41695 610
rect 41491 572 41537 582
rect 41621 572 41667 582
rect 41747 217 41817 713
rect 42149 679 42175 713
rect 41983 661 41994 672
rect 41943 611 41959 645
rect 41983 611 42015 661
rect 42125 651 42175 679
rect 42125 645 42141 651
rect 42143 611 42175 651
rect 41983 601 42017 611
rect 42141 601 42175 611
rect 41863 600 41965 601
rect 41983 600 42175 601
rect 41891 572 41937 573
rect 41983 319 42017 600
rect 42027 573 42051 577
rect 42107 573 42131 577
rect 42021 572 42067 573
rect 42027 353 42051 572
rect 42059 369 42061 561
rect 42063 400 42067 572
rect 42085 572 42137 573
rect 42085 357 42131 572
rect 42107 353 42131 357
rect 42141 353 42175 600
rect 42125 319 42175 353
rect 41943 285 41959 319
rect 41983 269 42015 319
rect 42143 269 42175 319
rect 41983 258 41994 269
rect 42149 217 42175 269
rect 42183 661 42217 713
rect 42349 679 42375 713
rect 42183 611 42215 661
rect 42325 651 42375 679
rect 42325 645 42341 651
rect 42343 611 42375 651
rect 42183 601 42217 611
rect 42341 601 42375 611
rect 42183 600 42375 601
rect 42183 319 42217 600
rect 42227 573 42251 577
rect 42307 573 42331 577
rect 42221 572 42267 573
rect 42227 353 42251 572
rect 42259 369 42261 561
rect 42263 400 42267 572
rect 42285 572 42337 573
rect 42285 357 42331 572
rect 42307 353 42331 357
rect 42341 353 42375 600
rect 42325 319 42375 353
rect 42183 269 42215 319
rect 42343 269 42375 319
rect 42183 217 42217 269
rect 42349 217 42375 269
rect 42383 661 42417 713
rect 42549 679 42575 713
rect 42383 611 42415 661
rect 42525 651 42575 679
rect 42525 645 42541 651
rect 42543 611 42575 651
rect 42383 601 42417 611
rect 42541 601 42575 611
rect 42383 600 42575 601
rect 42383 319 42417 600
rect 42427 573 42451 577
rect 42507 573 42531 577
rect 42421 572 42467 573
rect 42427 353 42451 572
rect 42459 369 42461 561
rect 42463 400 42467 572
rect 42485 572 42537 573
rect 42485 357 42531 572
rect 42507 353 42531 357
rect 42541 353 42575 600
rect 42525 319 42575 353
rect 42383 269 42415 319
rect 42543 269 42575 319
rect 42383 217 42417 269
rect 42549 217 42575 269
rect 42583 661 42617 713
rect 42749 679 42775 713
rect 42583 611 42615 661
rect 42725 651 42775 679
rect 42725 645 42741 651
rect 42743 611 42775 651
rect 42583 601 42617 611
rect 42741 601 42775 611
rect 42583 600 42775 601
rect 42583 319 42617 600
rect 42627 573 42651 577
rect 42707 573 42731 577
rect 42621 572 42667 573
rect 42627 353 42651 572
rect 42659 369 42661 561
rect 42663 400 42667 572
rect 42685 572 42737 573
rect 42685 357 42731 572
rect 42707 353 42731 357
rect 42741 353 42775 600
rect 42725 319 42775 353
rect 42583 269 42615 319
rect 42743 269 42775 319
rect 42583 217 42617 269
rect 42749 217 42775 269
rect 42783 661 42817 713
rect 42783 611 42815 661
rect 42925 651 42975 679
rect 42925 645 42941 651
rect 42943 611 42975 651
rect 42999 611 43009 645
rect 42783 601 42817 611
rect 42941 601 42975 611
rect 42783 600 42975 601
rect 42993 600 43095 601
rect 42783 319 42817 600
rect 42827 573 42851 577
rect 42907 573 42931 577
rect 42821 572 42867 573
rect 42827 353 42851 572
rect 42859 369 42861 561
rect 42863 400 42867 572
rect 42885 572 42937 573
rect 42885 357 42931 572
rect 42907 353 42931 357
rect 42941 353 42975 600
rect 43021 572 43067 573
rect 42925 319 42975 353
rect 42783 269 42815 319
rect 42943 269 42975 319
rect 42999 285 43009 319
rect 42783 217 42817 269
rect 42964 258 42975 269
rect 43147 217 43217 731
rect 43547 713 43629 747
rect 43679 713 44879 747
rect 44947 731 45029 749
rect 45329 747 45412 749
rect 46747 765 46811 783
rect 47147 765 47212 783
rect 46747 749 47212 765
rect 43263 600 43365 610
rect 43393 600 43495 610
rect 43291 572 43337 582
rect 43421 572 43467 582
rect 43547 217 43617 713
rect 43949 679 43975 713
rect 43783 661 43794 672
rect 43743 611 43759 645
rect 43783 611 43815 661
rect 43925 651 43975 679
rect 43925 645 43941 651
rect 43943 611 43975 651
rect 43783 601 43817 611
rect 43941 601 43975 611
rect 43663 600 43765 601
rect 43783 600 43975 601
rect 43691 572 43737 573
rect 43783 319 43817 600
rect 43827 573 43851 577
rect 43907 573 43931 577
rect 43821 572 43867 573
rect 43827 353 43851 572
rect 43859 369 43861 561
rect 43863 400 43867 572
rect 43885 572 43937 573
rect 43885 357 43931 572
rect 43907 353 43931 357
rect 43941 353 43975 600
rect 43925 319 43975 353
rect 43743 285 43759 319
rect 43783 269 43815 319
rect 43943 269 43975 319
rect 43783 258 43794 269
rect 43949 217 43975 269
rect 43983 661 44017 713
rect 44149 679 44175 713
rect 43983 611 44015 661
rect 44125 651 44175 679
rect 44125 645 44141 651
rect 44143 611 44175 651
rect 43983 601 44017 611
rect 44141 601 44175 611
rect 43983 600 44175 601
rect 43983 319 44017 600
rect 44027 573 44051 577
rect 44107 573 44131 577
rect 44021 572 44067 573
rect 44027 353 44051 572
rect 44059 369 44061 561
rect 44063 400 44067 572
rect 44085 572 44137 573
rect 44085 357 44131 572
rect 44107 353 44131 357
rect 44141 353 44175 600
rect 44125 319 44175 353
rect 43983 269 44015 319
rect 44143 269 44175 319
rect 43983 217 44017 269
rect 44149 217 44175 269
rect 44183 661 44217 713
rect 44349 679 44375 713
rect 44183 611 44215 661
rect 44325 651 44375 679
rect 44325 645 44341 651
rect 44343 611 44375 651
rect 44183 601 44217 611
rect 44341 601 44375 611
rect 44183 600 44375 601
rect 44183 319 44217 600
rect 44227 573 44251 577
rect 44307 573 44331 577
rect 44221 572 44267 573
rect 44227 353 44251 572
rect 44259 369 44261 561
rect 44263 400 44267 572
rect 44285 572 44337 573
rect 44285 357 44331 572
rect 44307 353 44331 357
rect 44341 353 44375 600
rect 44325 319 44375 353
rect 44183 269 44215 319
rect 44343 269 44375 319
rect 44183 217 44217 269
rect 44349 217 44375 269
rect 44383 661 44417 713
rect 44549 679 44575 713
rect 44383 611 44415 661
rect 44525 651 44575 679
rect 44525 645 44541 651
rect 44543 611 44575 651
rect 44383 601 44417 611
rect 44541 601 44575 611
rect 44383 600 44575 601
rect 44383 319 44417 600
rect 44427 573 44451 577
rect 44507 573 44531 577
rect 44421 572 44467 573
rect 44427 353 44451 572
rect 44459 369 44461 561
rect 44463 400 44467 572
rect 44485 572 44537 573
rect 44485 357 44531 572
rect 44507 353 44531 357
rect 44541 353 44575 600
rect 44525 319 44575 353
rect 44383 269 44415 319
rect 44543 269 44575 319
rect 44383 217 44417 269
rect 44549 217 44575 269
rect 44583 661 44617 713
rect 44583 611 44615 661
rect 44725 651 44775 679
rect 44725 645 44741 651
rect 44743 611 44775 651
rect 44799 611 44809 645
rect 44583 601 44617 611
rect 44741 601 44775 611
rect 44583 600 44775 601
rect 44793 600 44895 601
rect 44583 319 44617 600
rect 44627 573 44651 577
rect 44707 573 44731 577
rect 44621 572 44667 573
rect 44627 353 44651 572
rect 44659 369 44661 561
rect 44663 400 44667 572
rect 44685 572 44737 573
rect 44685 357 44731 572
rect 44707 353 44731 357
rect 44741 353 44775 600
rect 44821 572 44867 573
rect 44725 319 44775 353
rect 44583 269 44615 319
rect 44743 269 44775 319
rect 44799 285 44809 319
rect 44583 217 44617 269
rect 44764 258 44775 269
rect 44947 217 45017 731
rect 45347 713 45429 747
rect 45479 713 46679 747
rect 46747 731 46829 749
rect 47129 747 47212 749
rect 48547 765 48611 783
rect 48947 765 49012 783
rect 48547 749 49012 765
rect 45063 600 45165 610
rect 45193 600 45295 610
rect 45091 572 45137 582
rect 45221 572 45267 582
rect 45347 217 45417 713
rect 45749 679 45775 713
rect 45583 661 45594 672
rect 45543 611 45559 645
rect 45583 611 45615 661
rect 45725 651 45775 679
rect 45725 645 45741 651
rect 45743 611 45775 651
rect 45583 601 45617 611
rect 45741 601 45775 611
rect 45463 600 45565 601
rect 45583 600 45775 601
rect 45491 572 45537 573
rect 45583 319 45617 600
rect 45627 573 45651 577
rect 45707 573 45731 577
rect 45621 572 45667 573
rect 45627 353 45651 572
rect 45659 369 45661 561
rect 45663 400 45667 572
rect 45685 572 45737 573
rect 45685 357 45731 572
rect 45707 353 45731 357
rect 45741 353 45775 600
rect 45725 319 45775 353
rect 45543 285 45559 319
rect 45583 269 45615 319
rect 45743 269 45775 319
rect 45583 258 45594 269
rect 45749 217 45775 269
rect 45783 661 45817 713
rect 45949 679 45975 713
rect 45783 611 45815 661
rect 45925 651 45975 679
rect 45925 645 45941 651
rect 45943 611 45975 651
rect 45783 601 45817 611
rect 45941 601 45975 611
rect 45783 600 45975 601
rect 45783 319 45817 600
rect 45827 573 45851 577
rect 45907 573 45931 577
rect 45821 572 45867 573
rect 45827 353 45851 572
rect 45859 369 45861 561
rect 45863 400 45867 572
rect 45885 572 45937 573
rect 45885 357 45931 572
rect 45907 353 45931 357
rect 45941 353 45975 600
rect 45925 319 45975 353
rect 45783 269 45815 319
rect 45943 269 45975 319
rect 45783 217 45817 269
rect 45949 217 45975 269
rect 45983 661 46017 713
rect 46149 679 46175 713
rect 45983 611 46015 661
rect 46125 651 46175 679
rect 46125 645 46141 651
rect 46143 611 46175 651
rect 45983 601 46017 611
rect 46141 601 46175 611
rect 45983 600 46175 601
rect 45983 319 46017 600
rect 46027 573 46051 577
rect 46107 573 46131 577
rect 46021 572 46067 573
rect 46027 353 46051 572
rect 46059 369 46061 561
rect 46063 400 46067 572
rect 46085 572 46137 573
rect 46085 357 46131 572
rect 46107 353 46131 357
rect 46141 353 46175 600
rect 46125 319 46175 353
rect 45983 269 46015 319
rect 46143 269 46175 319
rect 45983 217 46017 269
rect 46149 217 46175 269
rect 46183 661 46217 713
rect 46349 679 46375 713
rect 46183 611 46215 661
rect 46325 651 46375 679
rect 46325 645 46341 651
rect 46343 611 46375 651
rect 46183 601 46217 611
rect 46341 601 46375 611
rect 46183 600 46375 601
rect 46183 319 46217 600
rect 46227 573 46251 577
rect 46307 573 46331 577
rect 46221 572 46267 573
rect 46227 353 46251 572
rect 46259 369 46261 561
rect 46263 400 46267 572
rect 46285 572 46337 573
rect 46285 357 46331 572
rect 46307 353 46331 357
rect 46341 353 46375 600
rect 46325 319 46375 353
rect 46183 269 46215 319
rect 46343 269 46375 319
rect 46183 217 46217 269
rect 46349 217 46375 269
rect 46383 661 46417 713
rect 46383 611 46415 661
rect 46525 651 46575 679
rect 46525 645 46541 651
rect 46543 611 46575 651
rect 46599 611 46609 645
rect 46383 601 46417 611
rect 46541 601 46575 611
rect 46383 600 46575 601
rect 46593 600 46695 601
rect 46383 319 46417 600
rect 46427 573 46451 577
rect 46507 573 46531 577
rect 46421 572 46467 573
rect 46427 353 46451 572
rect 46459 369 46461 561
rect 46463 400 46467 572
rect 46485 572 46537 573
rect 46485 357 46531 572
rect 46507 353 46531 357
rect 46541 353 46575 600
rect 46621 572 46667 573
rect 46525 319 46575 353
rect 46383 269 46415 319
rect 46543 269 46575 319
rect 46599 285 46609 319
rect 46383 217 46417 269
rect 46564 258 46575 269
rect 46747 217 46817 731
rect 47147 713 47229 747
rect 47279 713 48479 747
rect 48547 731 48629 749
rect 48929 747 49012 749
rect 50347 765 50411 783
rect 50747 765 50812 783
rect 50347 749 50812 765
rect 46863 600 46965 610
rect 46993 600 47095 610
rect 46891 572 46937 582
rect 47021 572 47067 582
rect 47147 217 47217 713
rect 47549 679 47575 713
rect 47383 661 47394 672
rect 47343 611 47359 645
rect 47383 611 47415 661
rect 47525 651 47575 679
rect 47525 645 47541 651
rect 47543 611 47575 651
rect 47383 601 47417 611
rect 47541 601 47575 611
rect 47263 600 47365 601
rect 47383 600 47575 601
rect 47291 572 47337 573
rect 47383 319 47417 600
rect 47427 573 47451 577
rect 47507 573 47531 577
rect 47421 572 47467 573
rect 47427 353 47451 572
rect 47459 369 47461 561
rect 47463 400 47467 572
rect 47485 572 47537 573
rect 47485 357 47531 572
rect 47507 353 47531 357
rect 47541 353 47575 600
rect 47525 319 47575 353
rect 47343 285 47359 319
rect 47383 269 47415 319
rect 47543 269 47575 319
rect 47383 258 47394 269
rect 47549 217 47575 269
rect 47583 661 47617 713
rect 47749 679 47775 713
rect 47583 611 47615 661
rect 47725 651 47775 679
rect 47725 645 47741 651
rect 47743 611 47775 651
rect 47583 601 47617 611
rect 47741 601 47775 611
rect 47583 600 47775 601
rect 47583 319 47617 600
rect 47627 573 47651 577
rect 47707 573 47731 577
rect 47621 572 47667 573
rect 47627 353 47651 572
rect 47659 369 47661 561
rect 47663 400 47667 572
rect 47685 572 47737 573
rect 47685 357 47731 572
rect 47707 353 47731 357
rect 47741 353 47775 600
rect 47725 319 47775 353
rect 47583 269 47615 319
rect 47743 269 47775 319
rect 47583 217 47617 269
rect 47749 217 47775 269
rect 47783 661 47817 713
rect 47949 679 47975 713
rect 47783 611 47815 661
rect 47925 651 47975 679
rect 47925 645 47941 651
rect 47943 611 47975 651
rect 47783 601 47817 611
rect 47941 601 47975 611
rect 47783 600 47975 601
rect 47783 319 47817 600
rect 47827 573 47851 577
rect 47907 573 47931 577
rect 47821 572 47867 573
rect 47827 353 47851 572
rect 47859 369 47861 561
rect 47863 400 47867 572
rect 47885 572 47937 573
rect 47885 357 47931 572
rect 47907 353 47931 357
rect 47941 353 47975 600
rect 47925 319 47975 353
rect 47783 269 47815 319
rect 47943 269 47975 319
rect 47783 217 47817 269
rect 47949 217 47975 269
rect 47983 661 48017 713
rect 48149 679 48175 713
rect 47983 611 48015 661
rect 48125 651 48175 679
rect 48125 645 48141 651
rect 48143 611 48175 651
rect 47983 601 48017 611
rect 48141 601 48175 611
rect 47983 600 48175 601
rect 47983 319 48017 600
rect 48027 573 48051 577
rect 48107 573 48131 577
rect 48021 572 48067 573
rect 48027 353 48051 572
rect 48059 369 48061 561
rect 48063 400 48067 572
rect 48085 572 48137 573
rect 48085 357 48131 572
rect 48107 353 48131 357
rect 48141 353 48175 600
rect 48125 319 48175 353
rect 47983 269 48015 319
rect 48143 269 48175 319
rect 47983 217 48017 269
rect 48149 217 48175 269
rect 48183 661 48217 713
rect 48183 611 48215 661
rect 48325 651 48375 679
rect 48325 645 48341 651
rect 48343 611 48375 651
rect 48399 611 48409 645
rect 48183 601 48217 611
rect 48341 601 48375 611
rect 48183 600 48375 601
rect 48393 600 48495 601
rect 48183 319 48217 600
rect 48227 573 48251 577
rect 48307 573 48331 577
rect 48221 572 48267 573
rect 48227 353 48251 572
rect 48259 369 48261 561
rect 48263 400 48267 572
rect 48285 572 48337 573
rect 48285 357 48331 572
rect 48307 353 48331 357
rect 48341 353 48375 600
rect 48421 572 48467 573
rect 48325 319 48375 353
rect 48183 269 48215 319
rect 48343 269 48375 319
rect 48399 285 48409 319
rect 48183 217 48217 269
rect 48364 258 48375 269
rect 48547 217 48617 731
rect 48947 713 49029 747
rect 49079 713 50279 747
rect 50347 731 50429 749
rect 50729 747 50812 749
rect 52147 765 52211 783
rect 52547 765 52612 783
rect 52147 749 52612 765
rect 48663 600 48765 610
rect 48793 600 48895 610
rect 48691 572 48737 582
rect 48821 572 48867 582
rect 48947 217 49017 713
rect 49349 679 49375 713
rect 49183 661 49194 672
rect 49143 611 49159 645
rect 49183 611 49215 661
rect 49325 651 49375 679
rect 49325 645 49341 651
rect 49343 611 49375 651
rect 49183 601 49217 611
rect 49341 601 49375 611
rect 49063 600 49165 601
rect 49183 600 49375 601
rect 49091 572 49137 573
rect 49183 319 49217 600
rect 49227 573 49251 577
rect 49307 573 49331 577
rect 49221 572 49267 573
rect 49227 353 49251 572
rect 49259 369 49261 561
rect 49263 400 49267 572
rect 49285 572 49337 573
rect 49285 357 49331 572
rect 49307 353 49331 357
rect 49341 353 49375 600
rect 49325 319 49375 353
rect 49143 285 49159 319
rect 49183 269 49215 319
rect 49343 269 49375 319
rect 49183 258 49194 269
rect 49349 217 49375 269
rect 49383 661 49417 713
rect 49549 679 49575 713
rect 49383 611 49415 661
rect 49525 651 49575 679
rect 49525 645 49541 651
rect 49543 611 49575 651
rect 49383 601 49417 611
rect 49541 601 49575 611
rect 49383 600 49575 601
rect 49383 319 49417 600
rect 49427 573 49451 577
rect 49507 573 49531 577
rect 49421 572 49467 573
rect 49427 353 49451 572
rect 49459 369 49461 561
rect 49463 400 49467 572
rect 49485 572 49537 573
rect 49485 357 49531 572
rect 49507 353 49531 357
rect 49541 353 49575 600
rect 49525 319 49575 353
rect 49383 269 49415 319
rect 49543 269 49575 319
rect 49383 217 49417 269
rect 49549 217 49575 269
rect 49583 661 49617 713
rect 49749 679 49775 713
rect 49583 611 49615 661
rect 49725 651 49775 679
rect 49725 645 49741 651
rect 49743 611 49775 651
rect 49583 601 49617 611
rect 49741 601 49775 611
rect 49583 600 49775 601
rect 49583 319 49617 600
rect 49627 573 49651 577
rect 49707 573 49731 577
rect 49621 572 49667 573
rect 49627 353 49651 572
rect 49659 369 49661 561
rect 49663 400 49667 572
rect 49685 572 49737 573
rect 49685 357 49731 572
rect 49707 353 49731 357
rect 49741 353 49775 600
rect 49725 319 49775 353
rect 49583 269 49615 319
rect 49743 269 49775 319
rect 49583 217 49617 269
rect 49749 217 49775 269
rect 49783 661 49817 713
rect 49949 679 49975 713
rect 49783 611 49815 661
rect 49925 651 49975 679
rect 49925 645 49941 651
rect 49943 611 49975 651
rect 49783 601 49817 611
rect 49941 601 49975 611
rect 49783 600 49975 601
rect 49783 319 49817 600
rect 49827 573 49851 577
rect 49907 573 49931 577
rect 49821 572 49867 573
rect 49827 353 49851 572
rect 49859 369 49861 561
rect 49863 400 49867 572
rect 49885 572 49937 573
rect 49885 357 49931 572
rect 49907 353 49931 357
rect 49941 353 49975 600
rect 49925 319 49975 353
rect 49783 269 49815 319
rect 49943 269 49975 319
rect 49783 217 49817 269
rect 49949 217 49975 269
rect 49983 661 50017 713
rect 49983 611 50015 661
rect 50125 651 50175 679
rect 50125 645 50141 651
rect 50143 611 50175 651
rect 50199 611 50209 645
rect 49983 601 50017 611
rect 50141 601 50175 611
rect 49983 600 50175 601
rect 50193 600 50295 601
rect 49983 319 50017 600
rect 50027 573 50051 577
rect 50107 573 50131 577
rect 50021 572 50067 573
rect 50027 353 50051 572
rect 50059 369 50061 561
rect 50063 400 50067 572
rect 50085 572 50137 573
rect 50085 357 50131 572
rect 50107 353 50131 357
rect 50141 353 50175 600
rect 50221 572 50267 573
rect 50125 319 50175 353
rect 49983 269 50015 319
rect 50143 269 50175 319
rect 50199 285 50209 319
rect 49983 217 50017 269
rect 50164 258 50175 269
rect 50347 217 50417 731
rect 50747 713 50829 747
rect 50879 713 52079 747
rect 52147 731 52229 749
rect 52529 747 52612 749
rect 53947 765 54011 783
rect 54347 765 54412 783
rect 53947 749 54412 765
rect 50463 600 50565 610
rect 50593 600 50695 610
rect 50491 572 50537 582
rect 50621 572 50667 582
rect 50747 217 50817 713
rect 51149 679 51175 713
rect 50983 661 50994 672
rect 50943 611 50959 645
rect 50983 611 51015 661
rect 51125 651 51175 679
rect 51125 645 51141 651
rect 51143 611 51175 651
rect 50983 601 51017 611
rect 51141 601 51175 611
rect 50863 600 50965 601
rect 50983 600 51175 601
rect 50891 572 50937 573
rect 50983 319 51017 600
rect 51027 573 51051 577
rect 51107 573 51131 577
rect 51021 572 51067 573
rect 51027 353 51051 572
rect 51059 369 51061 561
rect 51063 400 51067 572
rect 51085 572 51137 573
rect 51085 357 51131 572
rect 51107 353 51131 357
rect 51141 353 51175 600
rect 51125 319 51175 353
rect 50943 285 50959 319
rect 50983 269 51015 319
rect 51143 269 51175 319
rect 50983 258 50994 269
rect 51149 217 51175 269
rect 51183 661 51217 713
rect 51349 679 51375 713
rect 51183 611 51215 661
rect 51325 651 51375 679
rect 51325 645 51341 651
rect 51343 611 51375 651
rect 51183 601 51217 611
rect 51341 601 51375 611
rect 51183 600 51375 601
rect 51183 319 51217 600
rect 51227 573 51251 577
rect 51307 573 51331 577
rect 51221 572 51267 573
rect 51227 353 51251 572
rect 51259 369 51261 561
rect 51263 400 51267 572
rect 51285 572 51337 573
rect 51285 357 51331 572
rect 51307 353 51331 357
rect 51341 353 51375 600
rect 51325 319 51375 353
rect 51183 269 51215 319
rect 51343 269 51375 319
rect 51183 217 51217 269
rect 51349 217 51375 269
rect 51383 661 51417 713
rect 51549 679 51575 713
rect 51383 611 51415 661
rect 51525 651 51575 679
rect 51525 645 51541 651
rect 51543 611 51575 651
rect 51383 601 51417 611
rect 51541 601 51575 611
rect 51383 600 51575 601
rect 51383 319 51417 600
rect 51427 573 51451 577
rect 51507 573 51531 577
rect 51421 572 51467 573
rect 51427 353 51451 572
rect 51459 369 51461 561
rect 51463 400 51467 572
rect 51485 572 51537 573
rect 51485 357 51531 572
rect 51507 353 51531 357
rect 51541 353 51575 600
rect 51525 319 51575 353
rect 51383 269 51415 319
rect 51543 269 51575 319
rect 51383 217 51417 269
rect 51549 217 51575 269
rect 51583 661 51617 713
rect 51749 679 51775 713
rect 51583 611 51615 661
rect 51725 651 51775 679
rect 51725 645 51741 651
rect 51743 611 51775 651
rect 51583 601 51617 611
rect 51741 601 51775 611
rect 51583 600 51775 601
rect 51583 319 51617 600
rect 51627 573 51651 577
rect 51707 573 51731 577
rect 51621 572 51667 573
rect 51627 353 51651 572
rect 51659 369 51661 561
rect 51663 400 51667 572
rect 51685 572 51737 573
rect 51685 357 51731 572
rect 51707 353 51731 357
rect 51741 353 51775 600
rect 51725 319 51775 353
rect 51583 269 51615 319
rect 51743 269 51775 319
rect 51583 217 51617 269
rect 51749 217 51775 269
rect 51783 661 51817 713
rect 51783 611 51815 661
rect 51925 651 51975 679
rect 51925 645 51941 651
rect 51943 611 51975 651
rect 51999 611 52009 645
rect 51783 601 51817 611
rect 51941 601 51975 611
rect 51783 600 51975 601
rect 51993 600 52095 601
rect 51783 319 51817 600
rect 51827 573 51851 577
rect 51907 573 51931 577
rect 51821 572 51867 573
rect 51827 353 51851 572
rect 51859 369 51861 561
rect 51863 400 51867 572
rect 51885 572 51937 573
rect 51885 357 51931 572
rect 51907 353 51931 357
rect 51941 353 51975 600
rect 52021 572 52067 573
rect 51925 319 51975 353
rect 51783 269 51815 319
rect 51943 269 51975 319
rect 51999 285 52009 319
rect 51783 217 51817 269
rect 51964 258 51975 269
rect 52147 217 52217 731
rect 52547 713 52629 747
rect 52679 713 53879 747
rect 53947 731 54029 749
rect 54329 747 54412 749
rect 55747 765 55811 783
rect 56147 765 56212 783
rect 55747 749 56212 765
rect 52263 600 52365 610
rect 52393 600 52495 610
rect 52291 572 52337 582
rect 52421 572 52467 582
rect 52547 217 52617 713
rect 52949 679 52975 713
rect 52783 661 52794 672
rect 52743 611 52759 645
rect 52783 611 52815 661
rect 52925 651 52975 679
rect 52925 645 52941 651
rect 52943 611 52975 651
rect 52783 601 52817 611
rect 52941 601 52975 611
rect 52663 600 52765 601
rect 52783 600 52975 601
rect 52691 572 52737 573
rect 52783 319 52817 600
rect 52827 573 52851 577
rect 52907 573 52931 577
rect 52821 572 52867 573
rect 52827 353 52851 572
rect 52859 369 52861 561
rect 52863 400 52867 572
rect 52885 572 52937 573
rect 52885 357 52931 572
rect 52907 353 52931 357
rect 52941 353 52975 600
rect 52925 319 52975 353
rect 52743 285 52759 319
rect 52783 269 52815 319
rect 52943 269 52975 319
rect 52783 258 52794 269
rect 52949 217 52975 269
rect 52983 661 53017 713
rect 53149 679 53175 713
rect 52983 611 53015 661
rect 53125 651 53175 679
rect 53125 645 53141 651
rect 53143 611 53175 651
rect 52983 601 53017 611
rect 53141 601 53175 611
rect 52983 600 53175 601
rect 52983 319 53017 600
rect 53027 573 53051 577
rect 53107 573 53131 577
rect 53021 572 53067 573
rect 53027 353 53051 572
rect 53059 369 53061 561
rect 53063 400 53067 572
rect 53085 572 53137 573
rect 53085 357 53131 572
rect 53107 353 53131 357
rect 53141 353 53175 600
rect 53125 319 53175 353
rect 52983 269 53015 319
rect 53143 269 53175 319
rect 52983 217 53017 269
rect 53149 217 53175 269
rect 53183 661 53217 713
rect 53349 679 53375 713
rect 53183 611 53215 661
rect 53325 651 53375 679
rect 53325 645 53341 651
rect 53343 611 53375 651
rect 53183 601 53217 611
rect 53341 601 53375 611
rect 53183 600 53375 601
rect 53183 319 53217 600
rect 53227 573 53251 577
rect 53307 573 53331 577
rect 53221 572 53267 573
rect 53227 353 53251 572
rect 53259 369 53261 561
rect 53263 400 53267 572
rect 53285 572 53337 573
rect 53285 357 53331 572
rect 53307 353 53331 357
rect 53341 353 53375 600
rect 53325 319 53375 353
rect 53183 269 53215 319
rect 53343 269 53375 319
rect 53183 217 53217 269
rect 53349 217 53375 269
rect 53383 661 53417 713
rect 53549 679 53575 713
rect 53383 611 53415 661
rect 53525 651 53575 679
rect 53525 645 53541 651
rect 53543 611 53575 651
rect 53383 601 53417 611
rect 53541 601 53575 611
rect 53383 600 53575 601
rect 53383 319 53417 600
rect 53427 573 53451 577
rect 53507 573 53531 577
rect 53421 572 53467 573
rect 53427 353 53451 572
rect 53459 369 53461 561
rect 53463 400 53467 572
rect 53485 572 53537 573
rect 53485 357 53531 572
rect 53507 353 53531 357
rect 53541 353 53575 600
rect 53525 319 53575 353
rect 53383 269 53415 319
rect 53543 269 53575 319
rect 53383 217 53417 269
rect 53549 217 53575 269
rect 53583 661 53617 713
rect 53583 611 53615 661
rect 53725 651 53775 679
rect 53725 645 53741 651
rect 53743 611 53775 651
rect 53799 611 53809 645
rect 53583 601 53617 611
rect 53741 601 53775 611
rect 53583 600 53775 601
rect 53793 600 53895 601
rect 53583 319 53617 600
rect 53627 573 53651 577
rect 53707 573 53731 577
rect 53621 572 53667 573
rect 53627 353 53651 572
rect 53659 369 53661 561
rect 53663 400 53667 572
rect 53685 572 53737 573
rect 53685 357 53731 572
rect 53707 353 53731 357
rect 53741 353 53775 600
rect 53821 572 53867 573
rect 53725 319 53775 353
rect 53583 269 53615 319
rect 53743 269 53775 319
rect 53799 285 53809 319
rect 53583 217 53617 269
rect 53764 258 53775 269
rect 53947 217 54017 731
rect 54347 713 54429 747
rect 54479 713 55679 747
rect 55747 731 55829 749
rect 56129 747 56212 749
rect 57547 765 57611 783
rect 57947 765 58012 783
rect 57547 749 58012 765
rect 54063 600 54165 610
rect 54193 600 54295 610
rect 54091 572 54137 582
rect 54221 572 54267 582
rect 54347 217 54417 713
rect 54749 679 54775 713
rect 54583 661 54594 672
rect 54543 611 54559 645
rect 54583 611 54615 661
rect 54725 651 54775 679
rect 54725 645 54741 651
rect 54743 611 54775 651
rect 54583 601 54617 611
rect 54741 601 54775 611
rect 54463 600 54565 601
rect 54583 600 54775 601
rect 54491 572 54537 573
rect 54583 319 54617 600
rect 54627 573 54651 577
rect 54707 573 54731 577
rect 54621 572 54667 573
rect 54627 353 54651 572
rect 54659 369 54661 561
rect 54663 400 54667 572
rect 54685 572 54737 573
rect 54685 357 54731 572
rect 54707 353 54731 357
rect 54741 353 54775 600
rect 54725 319 54775 353
rect 54543 285 54559 319
rect 54583 269 54615 319
rect 54743 269 54775 319
rect 54583 258 54594 269
rect 54749 217 54775 269
rect 54783 661 54817 713
rect 54949 679 54975 713
rect 54783 611 54815 661
rect 54925 651 54975 679
rect 54925 645 54941 651
rect 54943 611 54975 651
rect 54783 601 54817 611
rect 54941 601 54975 611
rect 54783 600 54975 601
rect 54783 319 54817 600
rect 54827 573 54851 577
rect 54907 573 54931 577
rect 54821 572 54867 573
rect 54827 353 54851 572
rect 54859 369 54861 561
rect 54863 400 54867 572
rect 54885 572 54937 573
rect 54885 357 54931 572
rect 54907 353 54931 357
rect 54941 353 54975 600
rect 54925 319 54975 353
rect 54783 269 54815 319
rect 54943 269 54975 319
rect 54783 217 54817 269
rect 54949 217 54975 269
rect 54983 661 55017 713
rect 55149 679 55175 713
rect 54983 611 55015 661
rect 55125 651 55175 679
rect 55125 645 55141 651
rect 55143 611 55175 651
rect 54983 601 55017 611
rect 55141 601 55175 611
rect 54983 600 55175 601
rect 54983 319 55017 600
rect 55027 573 55051 577
rect 55107 573 55131 577
rect 55021 572 55067 573
rect 55027 353 55051 572
rect 55059 369 55061 561
rect 55063 400 55067 572
rect 55085 572 55137 573
rect 55085 357 55131 572
rect 55107 353 55131 357
rect 55141 353 55175 600
rect 55125 319 55175 353
rect 54983 269 55015 319
rect 55143 269 55175 319
rect 54983 217 55017 269
rect 55149 217 55175 269
rect 55183 661 55217 713
rect 55349 679 55375 713
rect 55183 611 55215 661
rect 55325 651 55375 679
rect 55325 645 55341 651
rect 55343 611 55375 651
rect 55183 601 55217 611
rect 55341 601 55375 611
rect 55183 600 55375 601
rect 55183 319 55217 600
rect 55227 573 55251 577
rect 55307 573 55331 577
rect 55221 572 55267 573
rect 55227 353 55251 572
rect 55259 369 55261 561
rect 55263 400 55267 572
rect 55285 572 55337 573
rect 55285 357 55331 572
rect 55307 353 55331 357
rect 55341 353 55375 600
rect 55325 319 55375 353
rect 55183 269 55215 319
rect 55343 269 55375 319
rect 55183 217 55217 269
rect 55349 217 55375 269
rect 55383 661 55417 713
rect 55383 611 55415 661
rect 55525 651 55575 679
rect 55525 645 55541 651
rect 55543 611 55575 651
rect 55599 611 55609 645
rect 55383 601 55417 611
rect 55541 601 55575 611
rect 55383 600 55575 601
rect 55593 600 55695 601
rect 55383 319 55417 600
rect 55427 573 55451 577
rect 55507 573 55531 577
rect 55421 572 55467 573
rect 55427 353 55451 572
rect 55459 369 55461 561
rect 55463 400 55467 572
rect 55485 572 55537 573
rect 55485 357 55531 572
rect 55507 353 55531 357
rect 55541 353 55575 600
rect 55621 572 55667 573
rect 55525 319 55575 353
rect 55383 269 55415 319
rect 55543 269 55575 319
rect 55599 285 55609 319
rect 55383 217 55417 269
rect 55564 258 55575 269
rect 55747 217 55817 731
rect 56147 713 56229 747
rect 56279 713 57479 747
rect 57547 731 57629 749
rect 57929 747 58012 749
rect 59347 765 59411 783
rect 59747 765 59812 783
rect 59347 749 59812 765
rect 55863 600 55965 610
rect 55993 600 56095 610
rect 55891 572 55937 582
rect 56021 572 56067 582
rect 56147 217 56217 713
rect 56549 679 56575 713
rect 56383 661 56394 672
rect 56343 611 56359 645
rect 56383 611 56415 661
rect 56525 651 56575 679
rect 56525 645 56541 651
rect 56543 611 56575 651
rect 56383 601 56417 611
rect 56541 601 56575 611
rect 56263 600 56365 601
rect 56383 600 56575 601
rect 56291 572 56337 573
rect 56383 319 56417 600
rect 56427 573 56451 577
rect 56507 573 56531 577
rect 56421 572 56467 573
rect 56427 353 56451 572
rect 56459 369 56461 561
rect 56463 400 56467 572
rect 56485 572 56537 573
rect 56485 357 56531 572
rect 56507 353 56531 357
rect 56541 353 56575 600
rect 56525 319 56575 353
rect 56343 285 56359 319
rect 56383 269 56415 319
rect 56543 269 56575 319
rect 56383 258 56394 269
rect 56549 217 56575 269
rect 56583 661 56617 713
rect 56749 679 56775 713
rect 56583 611 56615 661
rect 56725 651 56775 679
rect 56725 645 56741 651
rect 56743 611 56775 651
rect 56583 601 56617 611
rect 56741 601 56775 611
rect 56583 600 56775 601
rect 56583 319 56617 600
rect 56627 573 56651 577
rect 56707 573 56731 577
rect 56621 572 56667 573
rect 56627 353 56651 572
rect 56659 369 56661 561
rect 56663 400 56667 572
rect 56685 572 56737 573
rect 56685 357 56731 572
rect 56707 353 56731 357
rect 56741 353 56775 600
rect 56725 319 56775 353
rect 56583 269 56615 319
rect 56743 269 56775 319
rect 56583 217 56617 269
rect 56749 217 56775 269
rect 56783 661 56817 713
rect 56949 679 56975 713
rect 56783 611 56815 661
rect 56925 651 56975 679
rect 56925 645 56941 651
rect 56943 611 56975 651
rect 56783 601 56817 611
rect 56941 601 56975 611
rect 56783 600 56975 601
rect 56783 319 56817 600
rect 56827 573 56851 577
rect 56907 573 56931 577
rect 56821 572 56867 573
rect 56827 353 56851 572
rect 56859 369 56861 561
rect 56863 400 56867 572
rect 56885 572 56937 573
rect 56885 357 56931 572
rect 56907 353 56931 357
rect 56941 353 56975 600
rect 56925 319 56975 353
rect 56783 269 56815 319
rect 56943 269 56975 319
rect 56783 217 56817 269
rect 56949 217 56975 269
rect 56983 661 57017 713
rect 57149 679 57175 713
rect 56983 611 57015 661
rect 57125 651 57175 679
rect 57125 645 57141 651
rect 57143 611 57175 651
rect 56983 601 57017 611
rect 57141 601 57175 611
rect 56983 600 57175 601
rect 56983 319 57017 600
rect 57027 573 57051 577
rect 57107 573 57131 577
rect 57021 572 57067 573
rect 57027 353 57051 572
rect 57059 369 57061 561
rect 57063 400 57067 572
rect 57085 572 57137 573
rect 57085 357 57131 572
rect 57107 353 57131 357
rect 57141 353 57175 600
rect 57125 319 57175 353
rect 56983 269 57015 319
rect 57143 269 57175 319
rect 56983 217 57017 269
rect 57149 217 57175 269
rect 57183 661 57217 713
rect 57183 611 57215 661
rect 57325 651 57375 679
rect 57325 645 57341 651
rect 57343 611 57375 651
rect 57399 611 57409 645
rect 57183 601 57217 611
rect 57341 601 57375 611
rect 57183 600 57375 601
rect 57393 600 57495 601
rect 57183 319 57217 600
rect 57227 573 57251 577
rect 57307 573 57331 577
rect 57221 572 57267 573
rect 57227 353 57251 572
rect 57259 369 57261 561
rect 57263 400 57267 572
rect 57285 572 57337 573
rect 57285 357 57331 572
rect 57307 353 57331 357
rect 57341 353 57375 600
rect 57421 572 57467 573
rect 57325 319 57375 353
rect 57183 269 57215 319
rect 57343 269 57375 319
rect 57399 285 57409 319
rect 57183 217 57217 269
rect 57364 258 57375 269
rect 57547 217 57617 731
rect 57947 713 58029 747
rect 58079 713 59279 747
rect 59347 731 59429 749
rect 59729 747 59812 749
rect 61147 765 61211 783
rect 61547 765 61612 783
rect 61147 749 61612 765
rect 57663 600 57765 610
rect 57793 600 57895 610
rect 57691 572 57737 582
rect 57821 572 57867 582
rect 57947 217 58017 713
rect 58349 679 58375 713
rect 58183 661 58194 672
rect 58143 611 58159 645
rect 58183 611 58215 661
rect 58325 651 58375 679
rect 58325 645 58341 651
rect 58343 611 58375 651
rect 58183 601 58217 611
rect 58341 601 58375 611
rect 58063 600 58165 601
rect 58183 600 58375 601
rect 58091 572 58137 573
rect 58183 319 58217 600
rect 58227 573 58251 577
rect 58307 573 58331 577
rect 58221 572 58267 573
rect 58227 353 58251 572
rect 58259 369 58261 561
rect 58263 400 58267 572
rect 58285 572 58337 573
rect 58285 357 58331 572
rect 58307 353 58331 357
rect 58341 353 58375 600
rect 58325 319 58375 353
rect 58143 285 58159 319
rect 58183 269 58215 319
rect 58343 269 58375 319
rect 58183 258 58194 269
rect 58349 217 58375 269
rect 58383 661 58417 713
rect 58549 679 58575 713
rect 58383 611 58415 661
rect 58525 651 58575 679
rect 58525 645 58541 651
rect 58543 611 58575 651
rect 58383 601 58417 611
rect 58541 601 58575 611
rect 58383 600 58575 601
rect 58383 319 58417 600
rect 58427 573 58451 577
rect 58507 573 58531 577
rect 58421 572 58467 573
rect 58427 353 58451 572
rect 58459 369 58461 561
rect 58463 400 58467 572
rect 58485 572 58537 573
rect 58485 357 58531 572
rect 58507 353 58531 357
rect 58541 353 58575 600
rect 58525 319 58575 353
rect 58383 269 58415 319
rect 58543 269 58575 319
rect 58383 217 58417 269
rect 58549 217 58575 269
rect 58583 661 58617 713
rect 58749 679 58775 713
rect 58583 611 58615 661
rect 58725 651 58775 679
rect 58725 645 58741 651
rect 58743 611 58775 651
rect 58583 601 58617 611
rect 58741 601 58775 611
rect 58583 600 58775 601
rect 58583 319 58617 600
rect 58627 573 58651 577
rect 58707 573 58731 577
rect 58621 572 58667 573
rect 58627 353 58651 572
rect 58659 369 58661 561
rect 58663 400 58667 572
rect 58685 572 58737 573
rect 58685 357 58731 572
rect 58707 353 58731 357
rect 58741 353 58775 600
rect 58725 319 58775 353
rect 58583 269 58615 319
rect 58743 269 58775 319
rect 58583 217 58617 269
rect 58749 217 58775 269
rect 58783 661 58817 713
rect 58949 679 58975 713
rect 58783 611 58815 661
rect 58925 651 58975 679
rect 58925 645 58941 651
rect 58943 611 58975 651
rect 58783 601 58817 611
rect 58941 601 58975 611
rect 58783 600 58975 601
rect 58783 319 58817 600
rect 58827 573 58851 577
rect 58907 573 58931 577
rect 58821 572 58867 573
rect 58827 353 58851 572
rect 58859 369 58861 561
rect 58863 400 58867 572
rect 58885 572 58937 573
rect 58885 357 58931 572
rect 58907 353 58931 357
rect 58941 353 58975 600
rect 58925 319 58975 353
rect 58783 269 58815 319
rect 58943 269 58975 319
rect 58783 217 58817 269
rect 58949 217 58975 269
rect 58983 661 59017 713
rect 58983 611 59015 661
rect 59125 651 59175 679
rect 59125 645 59141 651
rect 59143 611 59175 651
rect 59199 611 59209 645
rect 58983 601 59017 611
rect 59141 601 59175 611
rect 58983 600 59175 601
rect 59193 600 59295 601
rect 58983 319 59017 600
rect 59027 573 59051 577
rect 59107 573 59131 577
rect 59021 572 59067 573
rect 59027 353 59051 572
rect 59059 369 59061 561
rect 59063 400 59067 572
rect 59085 572 59137 573
rect 59085 357 59131 572
rect 59107 353 59131 357
rect 59141 353 59175 600
rect 59221 572 59267 573
rect 59125 319 59175 353
rect 58983 269 59015 319
rect 59143 269 59175 319
rect 59199 285 59209 319
rect 58983 217 59017 269
rect 59164 258 59175 269
rect 59347 217 59417 731
rect 59747 713 59829 747
rect 59879 713 61079 747
rect 61147 731 61229 749
rect 61529 747 61612 749
rect 62947 765 63011 783
rect 63347 765 63412 783
rect 62947 749 63412 765
rect 59463 600 59565 610
rect 59593 600 59695 610
rect 59491 572 59537 582
rect 59621 572 59667 582
rect 59747 217 59817 713
rect 60149 679 60175 713
rect 59983 661 59994 672
rect 59943 611 59959 645
rect 59983 611 60015 661
rect 60125 651 60175 679
rect 60125 645 60141 651
rect 60143 611 60175 651
rect 59983 601 60017 611
rect 60141 601 60175 611
rect 59863 600 59965 601
rect 59983 600 60175 601
rect 59891 572 59937 573
rect 59983 319 60017 600
rect 60027 573 60051 577
rect 60107 573 60131 577
rect 60021 572 60067 573
rect 60027 353 60051 572
rect 60059 369 60061 561
rect 60063 400 60067 572
rect 60085 572 60137 573
rect 60085 357 60131 572
rect 60107 353 60131 357
rect 60141 353 60175 600
rect 60125 319 60175 353
rect 59943 285 59959 319
rect 59983 269 60015 319
rect 60143 269 60175 319
rect 59983 258 59994 269
rect 60149 217 60175 269
rect 60183 661 60217 713
rect 60349 679 60375 713
rect 60183 611 60215 661
rect 60325 651 60375 679
rect 60325 645 60341 651
rect 60343 611 60375 651
rect 60183 601 60217 611
rect 60341 601 60375 611
rect 60183 600 60375 601
rect 60183 319 60217 600
rect 60227 573 60251 577
rect 60307 573 60331 577
rect 60221 572 60267 573
rect 60227 353 60251 572
rect 60259 369 60261 561
rect 60263 400 60267 572
rect 60285 572 60337 573
rect 60285 357 60331 572
rect 60307 353 60331 357
rect 60341 353 60375 600
rect 60325 319 60375 353
rect 60183 269 60215 319
rect 60343 269 60375 319
rect 60183 217 60217 269
rect 60349 217 60375 269
rect 60383 661 60417 713
rect 60549 679 60575 713
rect 60383 611 60415 661
rect 60525 651 60575 679
rect 60525 645 60541 651
rect 60543 611 60575 651
rect 60383 601 60417 611
rect 60541 601 60575 611
rect 60383 600 60575 601
rect 60383 319 60417 600
rect 60427 573 60451 577
rect 60507 573 60531 577
rect 60421 572 60467 573
rect 60427 353 60451 572
rect 60459 369 60461 561
rect 60463 400 60467 572
rect 60485 572 60537 573
rect 60485 357 60531 572
rect 60507 353 60531 357
rect 60541 353 60575 600
rect 60525 319 60575 353
rect 60383 269 60415 319
rect 60543 269 60575 319
rect 60383 217 60417 269
rect 60549 217 60575 269
rect 60583 661 60617 713
rect 60749 679 60775 713
rect 60583 611 60615 661
rect 60725 651 60775 679
rect 60725 645 60741 651
rect 60743 611 60775 651
rect 60583 601 60617 611
rect 60741 601 60775 611
rect 60583 600 60775 601
rect 60583 319 60617 600
rect 60627 573 60651 577
rect 60707 573 60731 577
rect 60621 572 60667 573
rect 60627 353 60651 572
rect 60659 369 60661 561
rect 60663 400 60667 572
rect 60685 572 60737 573
rect 60685 357 60731 572
rect 60707 353 60731 357
rect 60741 353 60775 600
rect 60725 319 60775 353
rect 60583 269 60615 319
rect 60743 269 60775 319
rect 60583 217 60617 269
rect 60749 217 60775 269
rect 60783 661 60817 713
rect 60783 611 60815 661
rect 60925 651 60975 679
rect 60925 645 60941 651
rect 60943 611 60975 651
rect 60999 611 61009 645
rect 60783 601 60817 611
rect 60941 601 60975 611
rect 60783 600 60975 601
rect 60993 600 61095 601
rect 60783 319 60817 600
rect 60827 573 60851 577
rect 60907 573 60931 577
rect 60821 572 60867 573
rect 60827 353 60851 572
rect 60859 369 60861 561
rect 60863 400 60867 572
rect 60885 572 60937 573
rect 60885 357 60931 572
rect 60907 353 60931 357
rect 60941 353 60975 600
rect 61021 572 61067 573
rect 60925 319 60975 353
rect 60783 269 60815 319
rect 60943 269 60975 319
rect 60999 285 61009 319
rect 60783 217 60817 269
rect 60964 258 60975 269
rect 61147 217 61217 731
rect 61547 713 61629 747
rect 61679 713 62879 747
rect 62947 731 63029 749
rect 63329 747 63412 749
rect 64747 765 64811 783
rect 65147 765 65212 783
rect 64747 749 65212 765
rect 61263 600 61365 610
rect 61393 600 61495 610
rect 61291 572 61337 582
rect 61421 572 61467 582
rect 61547 217 61617 713
rect 61949 679 61975 713
rect 61783 661 61794 672
rect 61743 611 61759 645
rect 61783 611 61815 661
rect 61925 651 61975 679
rect 61925 645 61941 651
rect 61943 611 61975 651
rect 61783 601 61817 611
rect 61941 601 61975 611
rect 61663 600 61765 601
rect 61783 600 61975 601
rect 61691 572 61737 573
rect 61783 319 61817 600
rect 61827 573 61851 577
rect 61907 573 61931 577
rect 61821 572 61867 573
rect 61827 353 61851 572
rect 61859 369 61861 561
rect 61863 400 61867 572
rect 61885 572 61937 573
rect 61885 357 61931 572
rect 61907 353 61931 357
rect 61941 353 61975 600
rect 61925 319 61975 353
rect 61743 285 61759 319
rect 61783 269 61815 319
rect 61943 269 61975 319
rect 61783 258 61794 269
rect 61949 217 61975 269
rect 61983 661 62017 713
rect 62149 679 62175 713
rect 61983 611 62015 661
rect 62125 651 62175 679
rect 62125 645 62141 651
rect 62143 611 62175 651
rect 61983 601 62017 611
rect 62141 601 62175 611
rect 61983 600 62175 601
rect 61983 319 62017 600
rect 62027 573 62051 577
rect 62107 573 62131 577
rect 62021 572 62067 573
rect 62027 353 62051 572
rect 62059 369 62061 561
rect 62063 400 62067 572
rect 62085 572 62137 573
rect 62085 357 62131 572
rect 62107 353 62131 357
rect 62141 353 62175 600
rect 62125 319 62175 353
rect 61983 269 62015 319
rect 62143 269 62175 319
rect 61983 217 62017 269
rect 62149 217 62175 269
rect 62183 661 62217 713
rect 62349 679 62375 713
rect 62183 611 62215 661
rect 62325 651 62375 679
rect 62325 645 62341 651
rect 62343 611 62375 651
rect 62183 601 62217 611
rect 62341 601 62375 611
rect 62183 600 62375 601
rect 62183 319 62217 600
rect 62227 573 62251 577
rect 62307 573 62331 577
rect 62221 572 62267 573
rect 62227 353 62251 572
rect 62259 369 62261 561
rect 62263 400 62267 572
rect 62285 572 62337 573
rect 62285 357 62331 572
rect 62307 353 62331 357
rect 62341 353 62375 600
rect 62325 319 62375 353
rect 62183 269 62215 319
rect 62343 269 62375 319
rect 62183 217 62217 269
rect 62349 217 62375 269
rect 62383 661 62417 713
rect 62549 679 62575 713
rect 62383 611 62415 661
rect 62525 651 62575 679
rect 62525 645 62541 651
rect 62543 611 62575 651
rect 62383 601 62417 611
rect 62541 601 62575 611
rect 62383 600 62575 601
rect 62383 319 62417 600
rect 62427 573 62451 577
rect 62507 573 62531 577
rect 62421 572 62467 573
rect 62427 353 62451 572
rect 62459 369 62461 561
rect 62463 400 62467 572
rect 62485 572 62537 573
rect 62485 357 62531 572
rect 62507 353 62531 357
rect 62541 353 62575 600
rect 62525 319 62575 353
rect 62383 269 62415 319
rect 62543 269 62575 319
rect 62383 217 62417 269
rect 62549 217 62575 269
rect 62583 661 62617 713
rect 62583 611 62615 661
rect 62725 651 62775 679
rect 62725 645 62741 651
rect 62743 611 62775 651
rect 62799 611 62809 645
rect 62583 601 62617 611
rect 62741 601 62775 611
rect 62583 600 62775 601
rect 62793 600 62895 601
rect 62583 319 62617 600
rect 62627 573 62651 577
rect 62707 573 62731 577
rect 62621 572 62667 573
rect 62627 353 62651 572
rect 62659 369 62661 561
rect 62663 400 62667 572
rect 62685 572 62737 573
rect 62685 357 62731 572
rect 62707 353 62731 357
rect 62741 353 62775 600
rect 62821 572 62867 573
rect 62725 319 62775 353
rect 62583 269 62615 319
rect 62743 269 62775 319
rect 62799 285 62809 319
rect 62583 217 62617 269
rect 62764 258 62775 269
rect 62947 217 63017 731
rect 63347 713 63429 747
rect 63479 713 64679 747
rect 64747 731 64829 749
rect 65129 747 65212 749
rect 66547 765 66611 783
rect 66947 765 67012 783
rect 66547 749 67012 765
rect 63063 600 63165 610
rect 63193 600 63295 610
rect 63091 572 63137 582
rect 63221 572 63267 582
rect 63347 217 63417 713
rect 63749 679 63775 713
rect 63583 661 63594 672
rect 63543 611 63559 645
rect 63583 611 63615 661
rect 63725 651 63775 679
rect 63725 645 63741 651
rect 63743 611 63775 651
rect 63583 601 63617 611
rect 63741 601 63775 611
rect 63463 600 63565 601
rect 63583 600 63775 601
rect 63491 572 63537 573
rect 63583 319 63617 600
rect 63627 573 63651 577
rect 63707 573 63731 577
rect 63621 572 63667 573
rect 63627 353 63651 572
rect 63659 369 63661 561
rect 63663 400 63667 572
rect 63685 572 63737 573
rect 63685 357 63731 572
rect 63707 353 63731 357
rect 63741 353 63775 600
rect 63725 319 63775 353
rect 63543 285 63559 319
rect 63583 269 63615 319
rect 63743 269 63775 319
rect 63583 258 63594 269
rect 63749 217 63775 269
rect 63783 661 63817 713
rect 63949 679 63975 713
rect 63783 611 63815 661
rect 63925 651 63975 679
rect 63925 645 63941 651
rect 63943 611 63975 651
rect 63783 601 63817 611
rect 63941 601 63975 611
rect 63783 600 63975 601
rect 63783 319 63817 600
rect 63827 573 63851 577
rect 63907 573 63931 577
rect 63821 572 63867 573
rect 63827 353 63851 572
rect 63859 369 63861 561
rect 63863 400 63867 572
rect 63885 572 63937 573
rect 63885 357 63931 572
rect 63907 353 63931 357
rect 63941 353 63975 600
rect 63925 319 63975 353
rect 63783 269 63815 319
rect 63943 269 63975 319
rect 63783 217 63817 269
rect 63949 217 63975 269
rect 63983 661 64017 713
rect 64149 679 64175 713
rect 63983 611 64015 661
rect 64125 651 64175 679
rect 64125 645 64141 651
rect 64143 611 64175 651
rect 63983 601 64017 611
rect 64141 601 64175 611
rect 63983 600 64175 601
rect 63983 319 64017 600
rect 64027 573 64051 577
rect 64107 573 64131 577
rect 64021 572 64067 573
rect 64027 353 64051 572
rect 64059 369 64061 561
rect 64063 400 64067 572
rect 64085 572 64137 573
rect 64085 357 64131 572
rect 64107 353 64131 357
rect 64141 353 64175 600
rect 64125 319 64175 353
rect 63983 269 64015 319
rect 64143 269 64175 319
rect 63983 217 64017 269
rect 64149 217 64175 269
rect 64183 661 64217 713
rect 64349 679 64375 713
rect 64183 611 64215 661
rect 64325 651 64375 679
rect 64325 645 64341 651
rect 64343 611 64375 651
rect 64183 601 64217 611
rect 64341 601 64375 611
rect 64183 600 64375 601
rect 64183 319 64217 600
rect 64227 573 64251 577
rect 64307 573 64331 577
rect 64221 572 64267 573
rect 64227 353 64251 572
rect 64259 369 64261 561
rect 64263 400 64267 572
rect 64285 572 64337 573
rect 64285 357 64331 572
rect 64307 353 64331 357
rect 64341 353 64375 600
rect 64325 319 64375 353
rect 64183 269 64215 319
rect 64343 269 64375 319
rect 64183 217 64217 269
rect 64349 217 64375 269
rect 64383 661 64417 713
rect 64383 611 64415 661
rect 64525 651 64575 679
rect 64525 645 64541 651
rect 64543 611 64575 651
rect 64599 611 64609 645
rect 64383 601 64417 611
rect 64541 601 64575 611
rect 64383 600 64575 601
rect 64593 600 64695 601
rect 64383 319 64417 600
rect 64427 573 64451 577
rect 64507 573 64531 577
rect 64421 572 64467 573
rect 64427 353 64451 572
rect 64459 369 64461 561
rect 64463 400 64467 572
rect 64485 572 64537 573
rect 64485 357 64531 572
rect 64507 353 64531 357
rect 64541 353 64575 600
rect 64621 572 64667 573
rect 64525 319 64575 353
rect 64383 269 64415 319
rect 64543 269 64575 319
rect 64599 285 64609 319
rect 64383 217 64417 269
rect 64564 258 64575 269
rect 64747 217 64817 731
rect 65147 713 65229 747
rect 65279 713 66479 747
rect 66547 731 66629 749
rect 66929 747 67012 749
rect 68347 765 68411 783
rect 68347 749 68775 765
rect 64863 600 64965 610
rect 64993 600 65095 610
rect 64891 572 64937 582
rect 65021 572 65067 582
rect 65147 217 65217 713
rect 65549 679 65575 713
rect 65383 661 65394 672
rect 65343 611 65359 645
rect 65383 611 65415 661
rect 65525 651 65575 679
rect 65525 645 65541 651
rect 65543 611 65575 651
rect 65383 601 65417 611
rect 65541 601 65575 611
rect 65263 600 65365 601
rect 65383 600 65575 601
rect 65291 572 65337 573
rect 65383 319 65417 600
rect 65427 573 65451 577
rect 65507 573 65531 577
rect 65421 572 65467 573
rect 65427 353 65451 572
rect 65459 369 65461 561
rect 65463 400 65467 572
rect 65485 572 65537 573
rect 65485 357 65531 572
rect 65507 353 65531 357
rect 65541 353 65575 600
rect 65525 319 65575 353
rect 65343 285 65359 319
rect 65383 269 65415 319
rect 65543 269 65575 319
rect 65383 258 65394 269
rect 65549 217 65575 269
rect 65583 661 65617 713
rect 65749 679 65775 713
rect 65583 611 65615 661
rect 65725 651 65775 679
rect 65725 645 65741 651
rect 65743 611 65775 651
rect 65583 601 65617 611
rect 65741 601 65775 611
rect 65583 600 65775 601
rect 65583 319 65617 600
rect 65627 573 65651 577
rect 65707 573 65731 577
rect 65621 572 65667 573
rect 65627 353 65651 572
rect 65659 369 65661 561
rect 65663 400 65667 572
rect 65685 572 65737 573
rect 65685 357 65731 572
rect 65707 353 65731 357
rect 65741 353 65775 600
rect 65725 319 65775 353
rect 65583 269 65615 319
rect 65743 269 65775 319
rect 65583 217 65617 269
rect 65749 217 65775 269
rect 65783 661 65817 713
rect 65949 679 65975 713
rect 65783 611 65815 661
rect 65925 651 65975 679
rect 65925 645 65941 651
rect 65943 611 65975 651
rect 65783 601 65817 611
rect 65941 601 65975 611
rect 65783 600 65975 601
rect 65783 319 65817 600
rect 65827 573 65851 577
rect 65907 573 65931 577
rect 65821 572 65867 573
rect 65827 353 65851 572
rect 65859 369 65861 561
rect 65863 400 65867 572
rect 65885 572 65937 573
rect 65885 357 65931 572
rect 65907 353 65931 357
rect 65941 353 65975 600
rect 65925 319 65975 353
rect 65783 269 65815 319
rect 65943 269 65975 319
rect 65783 217 65817 269
rect 65949 217 65975 269
rect 65983 661 66017 713
rect 66149 679 66175 713
rect 65983 611 66015 661
rect 66125 651 66175 679
rect 66125 645 66141 651
rect 66143 611 66175 651
rect 65983 601 66017 611
rect 66141 601 66175 611
rect 65983 600 66175 601
rect 65983 319 66017 600
rect 66027 573 66051 577
rect 66107 573 66131 577
rect 66021 572 66067 573
rect 66027 353 66051 572
rect 66059 369 66061 561
rect 66063 400 66067 572
rect 66085 572 66137 573
rect 66085 357 66131 572
rect 66107 353 66131 357
rect 66141 353 66175 600
rect 66125 319 66175 353
rect 65983 269 66015 319
rect 66143 269 66175 319
rect 65983 217 66017 269
rect 66149 217 66175 269
rect 66183 661 66217 713
rect 66183 611 66215 661
rect 66325 651 66375 679
rect 66325 645 66341 651
rect 66343 611 66375 651
rect 66399 611 66409 645
rect 66183 601 66217 611
rect 66341 601 66375 611
rect 66183 600 66375 601
rect 66393 600 66495 601
rect 66183 319 66217 600
rect 66227 573 66251 577
rect 66307 573 66331 577
rect 66221 572 66267 573
rect 66227 353 66251 572
rect 66259 369 66261 561
rect 66263 400 66267 572
rect 66285 572 66337 573
rect 66285 357 66331 572
rect 66307 353 66331 357
rect 66341 353 66375 600
rect 66421 572 66467 573
rect 66325 319 66375 353
rect 66183 269 66215 319
rect 66343 269 66375 319
rect 66399 285 66409 319
rect 66183 217 66217 269
rect 66364 258 66375 269
rect 66547 217 66617 731
rect 66947 713 67029 747
rect 67079 713 68279 747
rect 68347 731 68429 749
rect 66663 600 66765 610
rect 66793 600 66895 610
rect 66691 572 66737 582
rect 66821 572 66867 582
rect 66947 217 67017 713
rect 67349 679 67375 713
rect 67183 661 67194 672
rect 67143 611 67159 645
rect 67183 611 67215 661
rect 67325 651 67375 679
rect 67325 645 67341 651
rect 67343 611 67375 651
rect 67183 601 67217 611
rect 67341 601 67375 611
rect 67063 600 67165 601
rect 67183 600 67375 601
rect 67091 572 67137 573
rect 67183 319 67217 600
rect 67227 573 67251 577
rect 67307 573 67331 577
rect 67221 572 67267 573
rect 67227 353 67251 572
rect 67259 369 67261 561
rect 67263 400 67267 572
rect 67285 572 67337 573
rect 67285 357 67331 572
rect 67307 353 67331 357
rect 67341 353 67375 600
rect 67325 319 67375 353
rect 67143 285 67159 319
rect 67183 269 67215 319
rect 67343 269 67375 319
rect 67183 258 67194 269
rect 67349 217 67375 269
rect 67383 661 67417 713
rect 67549 679 67575 713
rect 67383 611 67415 661
rect 67525 651 67575 679
rect 67525 645 67541 651
rect 67543 611 67575 651
rect 67383 601 67417 611
rect 67541 601 67575 611
rect 67383 600 67575 601
rect 67383 319 67417 600
rect 67427 573 67451 577
rect 67507 573 67531 577
rect 67421 572 67467 573
rect 67427 353 67451 572
rect 67459 369 67461 561
rect 67463 400 67467 572
rect 67485 572 67537 573
rect 67485 357 67531 572
rect 67507 353 67531 357
rect 67541 353 67575 600
rect 67525 319 67575 353
rect 67383 269 67415 319
rect 67543 269 67575 319
rect 67383 217 67417 269
rect 67549 217 67575 269
rect 67583 661 67617 713
rect 67749 679 67775 713
rect 67583 611 67615 661
rect 67725 651 67775 679
rect 67725 645 67741 651
rect 67743 611 67775 651
rect 67583 601 67617 611
rect 67741 601 67775 611
rect 67583 600 67775 601
rect 67583 319 67617 600
rect 67627 573 67651 577
rect 67707 573 67731 577
rect 67621 572 67667 573
rect 67627 353 67651 572
rect 67659 369 67661 561
rect 67663 400 67667 572
rect 67685 572 67737 573
rect 67685 357 67731 572
rect 67707 353 67731 357
rect 67741 353 67775 600
rect 67725 319 67775 353
rect 67583 269 67615 319
rect 67743 269 67775 319
rect 67583 217 67617 269
rect 67749 217 67775 269
rect 67783 661 67817 713
rect 67949 679 67975 713
rect 67783 611 67815 661
rect 67925 651 67975 679
rect 67925 645 67941 651
rect 67943 611 67975 651
rect 67783 601 67817 611
rect 67941 601 67975 611
rect 67783 600 67975 601
rect 67783 319 67817 600
rect 67827 573 67851 577
rect 67907 573 67931 577
rect 67821 572 67867 573
rect 67827 353 67851 572
rect 67859 369 67861 561
rect 67863 400 67867 572
rect 67885 572 67937 573
rect 67885 357 67931 572
rect 67907 353 67931 357
rect 67941 353 67975 600
rect 67925 319 67975 353
rect 67783 269 67815 319
rect 67943 269 67975 319
rect 67783 217 67817 269
rect 67949 217 67975 269
rect 67983 661 68017 713
rect 67983 611 68015 661
rect 68125 651 68175 679
rect 68125 645 68141 651
rect 68143 611 68175 651
rect 68199 611 68209 645
rect 67983 601 68017 611
rect 68141 601 68175 611
rect 67983 600 68175 601
rect 68193 600 68295 601
rect 67983 319 68017 600
rect 68027 573 68051 577
rect 68107 573 68131 577
rect 68021 572 68067 573
rect 68027 353 68051 572
rect 68059 369 68061 561
rect 68063 400 68067 572
rect 68085 572 68137 573
rect 68085 357 68131 572
rect 68107 353 68131 357
rect 68141 353 68175 600
rect 68221 572 68267 573
rect 68125 319 68175 353
rect 67983 269 68015 319
rect 68143 269 68175 319
rect 68199 285 68209 319
rect 67983 217 68017 269
rect 68164 258 68175 269
rect 68347 217 68417 731
rect 68463 600 68565 610
rect 68593 600 68695 610
rect 68491 572 68537 582
rect 68621 572 68667 582
rect 19783 183 19829 217
rect 20147 183 20229 217
rect 20279 183 21479 217
rect 21547 183 21629 217
rect 21947 183 22029 217
rect 22079 183 23279 217
rect 23347 183 23429 217
rect 23747 183 23829 217
rect 23879 183 25079 217
rect 25147 183 25229 217
rect 25547 183 25629 217
rect 25679 183 26879 217
rect 26947 183 27029 217
rect 27347 183 27429 217
rect 27479 183 28679 217
rect 28747 183 28829 217
rect 29147 183 29229 217
rect 29279 183 30479 217
rect 30547 183 30629 217
rect 30947 183 31029 217
rect 31079 183 32279 217
rect 32347 183 32429 217
rect 32747 183 32829 217
rect 32879 183 34079 217
rect 34147 183 34229 217
rect 34547 183 34629 217
rect 34679 183 35879 217
rect 35947 183 36029 217
rect 36347 183 36429 217
rect 36479 183 37679 217
rect 37747 183 37829 217
rect 38147 183 38229 217
rect 38279 183 39479 217
rect 39547 183 39629 217
rect 39947 183 40029 217
rect 40079 183 41279 217
rect 41347 183 41429 217
rect 41747 183 41829 217
rect 41879 183 43079 217
rect 43147 183 43229 217
rect 43547 183 43629 217
rect 43679 183 44879 217
rect 44947 183 45029 217
rect 45347 183 45429 217
rect 45479 183 46679 217
rect 46747 183 46829 217
rect 47147 183 47229 217
rect 47279 183 48479 217
rect 48547 183 48629 217
rect 48947 183 49029 217
rect 49079 183 50279 217
rect 50347 183 50429 217
rect 50747 183 50829 217
rect 50879 183 52079 217
rect 52147 183 52229 217
rect 52547 183 52629 217
rect 52679 183 53879 217
rect 53947 183 54029 217
rect 54347 183 54429 217
rect 54479 183 55679 217
rect 55747 183 55829 217
rect 56147 183 56229 217
rect 56279 183 57479 217
rect 57547 183 57629 217
rect 57947 183 58029 217
rect 58079 183 59279 217
rect 59347 183 59429 217
rect 59747 183 59829 217
rect 59879 183 61079 217
rect 61147 183 61229 217
rect 61547 183 61629 217
rect 61679 183 62879 217
rect 62947 183 63029 217
rect 63347 183 63429 217
rect 63479 183 64679 217
rect 64747 183 64829 217
rect 65147 183 65229 217
rect 65279 183 66479 217
rect 66547 183 66629 217
rect 66947 183 67029 217
rect 67079 183 68279 217
rect 68347 183 68429 217
rect 1147 147 1211 183
rect 3947 147 4011 183
rect 4747 147 4811 183
rect 8947 147 9011 183
rect 9347 147 9411 183
rect 10747 147 10811 183
rect 11147 147 11211 183
rect 12547 147 12611 183
rect 12947 147 13011 183
rect 14347 147 14411 183
rect 14747 147 14811 183
rect 16147 147 16211 183
rect 16547 147 16611 183
rect 19347 147 19411 183
rect 20147 147 20211 183
rect 21547 147 21611 183
rect 21947 147 22011 183
rect 23347 147 23411 183
rect 23747 147 23811 183
rect 25147 147 25211 183
rect 25547 147 25611 183
rect 26947 147 27011 183
rect 27347 147 27411 183
rect 28747 147 28811 183
rect 29147 147 29211 183
rect 30547 147 30611 183
rect 30947 147 31011 183
rect 32347 147 32411 183
rect 32747 147 32811 183
rect 34147 147 34211 183
rect 34547 147 34611 183
rect 35947 147 36011 183
rect 36347 147 36411 183
rect 37747 147 37811 183
rect 38147 147 38211 183
rect 39547 147 39611 183
rect 39947 147 40011 183
rect 41347 147 41411 183
rect 41747 147 41811 183
rect 43147 147 43211 183
rect 43547 147 43611 183
rect 44947 147 45011 183
rect 45347 147 45411 183
rect 46747 147 46811 183
rect 47147 147 47211 183
rect 48547 147 48611 183
rect 48947 147 49011 183
rect 50347 147 50411 183
rect 50747 147 50811 183
rect 52147 147 52211 183
rect 52547 147 52611 183
rect 53947 147 54011 183
rect 54347 147 54411 183
rect 55747 147 55811 183
rect 56147 147 56211 183
rect 57547 147 57611 183
rect 57947 147 58011 183
rect 59347 147 59411 183
rect 59747 147 59811 183
rect 61147 147 61211 183
rect 61547 147 61611 183
rect 62947 147 63011 183
rect 63347 147 63411 183
rect 64747 147 64811 183
rect 65147 147 65211 183
rect 66547 147 66611 183
rect 66947 147 67011 183
rect 68347 147 68411 183
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use SUNTR_NCHLCM  SUNTR_NCHLCM_0
timestamp 1713382353
transform 1 0 0 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_1
timestamp 1713382353
transform 1 0 809 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_2
timestamp 1713382353
transform 1 0 1015 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_3
timestamp 1713382353
transform 1 0 1623 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_4
timestamp 1713382353
transform 1 0 1829 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_5
timestamp 1713382353
transform 1 0 2035 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_6
timestamp 1713382353
transform 1 0 2442 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_7
timestamp 1713382353
transform 1 0 2849 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_8
timestamp 1713382353
transform 1 0 3256 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_9
timestamp 1713382353
transform 1 0 3663 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_10
timestamp 1713382353
transform 1 0 4070 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_11
timestamp 1713382353
transform 1 0 4276 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_12
timestamp 1713382353
transform 1 0 4884 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_13
timestamp 1713382353
transform 1 0 5291 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_14
timestamp 1713382353
transform 1 0 5698 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_15
timestamp 1713382353
transform 1 0 6105 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_16
timestamp 1713382353
transform 1 0 6512 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_17
timestamp 1713382353
transform 1 0 6919 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_18
timestamp 1713382353
transform 1 0 7326 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_19
timestamp 1713382353
transform 1 0 7733 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_20
timestamp 1713382353
transform 1 0 8140 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_21
timestamp 1713382353
transform 1 0 8547 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_22
timestamp 1713382353
transform 1 0 8954 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_23
timestamp 1713382353
transform 1 0 9361 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_24
timestamp 1713382353
transform 1 0 9768 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_25
timestamp 1713382353
transform 1 0 10175 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_26
timestamp 1713382353
transform 1 0 10582 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_27
timestamp 1713382353
transform 1 0 10989 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_28
timestamp 1713382353
transform 1 0 11396 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_29
timestamp 1713382353
transform 1 0 11803 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_30
timestamp 1713382353
transform 1 0 12210 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_31
timestamp 1713382353
transform 1 0 12617 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_32
timestamp 1713382353
transform 1 0 13024 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_33
timestamp 1713382353
transform 1 0 13431 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_34
timestamp 1713382353
transform 1 0 13838 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_35
timestamp 1713382353
transform 1 0 14245 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_36
timestamp 1713382353
transform 1 0 14652 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_37
timestamp 1713382353
transform 1 0 15059 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_38
timestamp 1713382353
transform 1 0 15466 0 1 1800
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_39
timestamp 1713382353
transform 1 0 1200 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_40
timestamp 1713382353
transform 1 0 2600 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_41
timestamp 1713382353
transform 1 0 4800 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_42
timestamp 1713382353
transform 1 0 6200 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_43
timestamp 1713382353
transform 1 0 7600 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_44
timestamp 1713382353
transform 1 0 9400 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_45
timestamp 1713382353
transform 1 0 11200 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_46
timestamp 1713382353
transform 1 0 13000 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_47
timestamp 1713382353
transform 1 0 14800 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_48
timestamp 1713382353
transform 1 0 16600 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_49
timestamp 1713382353
transform 1 0 18000 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_50
timestamp 1713382353
transform 1 0 20200 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_51
timestamp 1713382353
transform 1 0 22000 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_52
timestamp 1713382353
transform 1 0 23800 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_53
timestamp 1713382353
transform 1 0 25600 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_54
timestamp 1713382353
transform 1 0 27400 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_55
timestamp 1713382353
transform 1 0 29200 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_56
timestamp 1713382353
transform 1 0 31000 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_57
timestamp 1713382353
transform 1 0 32800 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_58
timestamp 1713382353
transform 1 0 34600 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_59
timestamp 1713382353
transform 1 0 36400 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_60
timestamp 1713382353
transform 1 0 38200 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_61
timestamp 1713382353
transform 1 0 40000 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_62
timestamp 1713382353
transform 1 0 41800 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_63
timestamp 1713382353
transform 1 0 43600 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_64
timestamp 1713382353
transform 1 0 45400 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_65
timestamp 1713382353
transform 1 0 47200 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_66
timestamp 1713382353
transform 1 0 49000 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_67
timestamp 1713382353
transform 1 0 50800 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_68
timestamp 1713382353
transform 1 0 52600 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_69
timestamp 1713382353
transform 1 0 54400 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_70
timestamp 1713382353
transform 1 0 56200 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_71
timestamp 1713382353
transform 1 0 58000 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_72
timestamp 1713382353
transform 1 0 59800 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_73
timestamp 1713382353
transform 1 0 61600 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_74
timestamp 1713382353
transform 1 0 63400 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_75
timestamp 1713382353
transform 1 0 65200 0 1 -400
box -53 -1200 1611 2983
use SUNTR_NCHLCM  SUNTR_NCHLCM_76
timestamp 1713382353
transform 1 0 67000 0 1 -400
box -53 -1200 1611 2983
use SUNTR_PCHLCM  SUNTR_PCHLCM_0
timestamp 1713382353
transform 1 0 206 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_1
timestamp 1713382353
transform 1 0 407 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_2
timestamp 1713382353
transform 1 0 608 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_3
timestamp 1713382353
transform 1 0 1221 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_4
timestamp 1713382353
transform 1 0 1422 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_5
timestamp 1713382353
transform 1 0 2241 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_6
timestamp 1713382353
transform 1 0 2648 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_7
timestamp 1713382353
transform 1 0 3055 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_8
timestamp 1713382353
transform 1 0 3462 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_9
timestamp 1713382353
transform 1 0 3869 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_10
timestamp 1713382353
transform 1 0 4482 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_11
timestamp 1713382353
transform 1 0 4683 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_12
timestamp 1713382353
transform 1 0 5090 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_13
timestamp 1713382353
transform 1 0 5497 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_14
timestamp 1713382353
transform 1 0 5904 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_15
timestamp 1713382353
transform 1 0 6311 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_16
timestamp 1713382353
transform 1 0 6718 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_17
timestamp 1713382353
transform 1 0 7125 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_18
timestamp 1713382353
transform 1 0 7532 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_19
timestamp 1713382353
transform 1 0 7939 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_20
timestamp 1713382353
transform 1 0 8346 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_21
timestamp 1713382353
transform 1 0 8753 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_22
timestamp 1713382353
transform 1 0 9160 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_23
timestamp 1713382353
transform 1 0 9567 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_24
timestamp 1713382353
transform 1 0 9974 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_25
timestamp 1713382353
transform 1 0 10381 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_26
timestamp 1713382353
transform 1 0 10788 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_27
timestamp 1713382353
transform 1 0 11195 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_28
timestamp 1713382353
transform 1 0 11602 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_29
timestamp 1713382353
transform 1 0 12009 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_30
timestamp 1713382353
transform 1 0 12416 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_31
timestamp 1713382353
transform 1 0 12823 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_32
timestamp 1713382353
transform 1 0 13230 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_33
timestamp 1713382353
transform 1 0 13637 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_34
timestamp 1713382353
transform 1 0 14044 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_35
timestamp 1713382353
transform 1 0 14451 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_36
timestamp 1713382353
transform 1 0 14858 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_37
timestamp 1713382353
transform 1 0 15265 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_38
timestamp 1713382353
transform 1 0 15672 0 1 1800
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_39
timestamp 1713382353
transform 1 0 0 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_40
timestamp 1713382353
transform 1 0 400 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_41
timestamp 1713382353
transform 1 0 800 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_42
timestamp 1713382353
transform 1 0 4000 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_43
timestamp 1713382353
transform 1 0 4400 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_44
timestamp 1713382353
transform 1 0 9000 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_45
timestamp 1713382353
transform 1 0 10800 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_46
timestamp 1713382353
transform 1 0 12600 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_47
timestamp 1713382353
transform 1 0 14400 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_48
timestamp 1713382353
transform 1 0 16200 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_49
timestamp 1713382353
transform 1 0 19400 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_50
timestamp 1713382353
transform 1 0 19800 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_51
timestamp 1713382353
transform 1 0 21600 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_52
timestamp 1713382353
transform 1 0 23400 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_53
timestamp 1713382353
transform 1 0 25200 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_54
timestamp 1713382353
transform 1 0 27000 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_55
timestamp 1713382353
transform 1 0 28800 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_56
timestamp 1713382353
transform 1 0 30600 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_57
timestamp 1713382353
transform 1 0 32400 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_58
timestamp 1713382353
transform 1 0 34200 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_59
timestamp 1713382353
transform 1 0 36000 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_60
timestamp 1713382353
transform 1 0 37800 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_61
timestamp 1713382353
transform 1 0 39600 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_62
timestamp 1713382353
transform 1 0 41400 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_63
timestamp 1713382353
transform 1 0 43200 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_64
timestamp 1713382353
transform 1 0 45000 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_65
timestamp 1713382353
transform 1 0 46800 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_66
timestamp 1713382353
transform 1 0 48600 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_67
timestamp 1713382353
transform 1 0 50400 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_68
timestamp 1713382353
transform 1 0 52200 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_69
timestamp 1713382353
transform 1 0 54000 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_70
timestamp 1713382353
transform 1 0 55800 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_71
timestamp 1713382353
transform 1 0 57600 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_72
timestamp 1713382353
transform 1 0 59400 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_73
timestamp 1713382353
transform 1 0 61200 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_74
timestamp 1713382353
transform 1 0 63000 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_75
timestamp 1713382353
transform 1 0 64800 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_76
timestamp 1713382353
transform 1 0 66600 0 1 -400
box -53 -1200 611 3001
use SUNTR_PCHLCM  SUNTR_PCHLCM_77
timestamp 1713382353
transform 1 0 68400 0 1 -400
box -53 -1200 611 3001
use SUNTR_NCHLCM  x1
timestamp 1713382353
transform 1 0 0 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x2
timestamp 1713382353
transform 1 0 2 0 1 600
box -53 -1200 611 3001
use SUNTR_PCHLCM  x3
timestamp 1713382353
transform 1 0 3 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x4
timestamp 1713382353
transform 1 0 4 0 1 600
box -53 -1200 1611 2983
use SUNTR_NCHLCM  x5
timestamp 1713382353
transform 1 0 5 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x6
timestamp 1713382353
transform 1 0 6 0 1 600
box -53 -1200 611 3001
use SUNTR_PCHLCM  x7
timestamp 1713382353
transform 1 0 7 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x8
timestamp 1713382353
transform 1 0 8 0 1 600
box -53 -1200 1611 2983
use SUNTR_NCHLCM  x9
timestamp 1713382353
transform 1 0 9 0 1 600
box -53 -1200 1611 2983
use SUNTR_NCHLCM  x10
timestamp 1713382353
transform 1 0 10 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x11
timestamp 1713382353
transform 1 0 11 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x12
timestamp 1713382353
transform 1 0 12 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x13
timestamp 1713382353
transform 1 0 13 0 1 600
box -53 -1200 611 3001
use SUNTR_PCHLCM  x14
timestamp 1713382353
transform 1 0 1 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x15
timestamp 1713382353
transform 1 0 14 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x16
timestamp 1713382353
transform 1 0 15 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x17
timestamp 1713382353
transform 1 0 16 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x18
timestamp 1713382353
transform 1 0 17 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x19
timestamp 1713382353
transform 1 0 18 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x20
timestamp 1713382353
transform 1 0 19 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x21
timestamp 1713382353
transform 1 0 20 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x22
timestamp 1713382353
transform 1 0 23 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x23
timestamp 1713382353
transform 1 0 24 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x24
timestamp 1713382353
transform 1 0 25 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x25
timestamp 1713382353
transform 1 0 21 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x26
timestamp 1713382353
transform 1 0 22 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x27
timestamp 1713382353
transform 1 0 26 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x28
timestamp 1713382353
transform 1 0 27 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x29
timestamp 1713382353
transform 1 0 28 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x30
timestamp 1713382353
transform 1 0 29 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x31
timestamp 1713382353
transform 1 0 30 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x32
timestamp 1713382353
transform 1 0 31 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x33
timestamp 1713382353
transform 1 0 32 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x34
timestamp 1713382353
transform 1 0 33 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x35
timestamp 1713382353
transform 1 0 34 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x36
timestamp 1713382353
transform 1 0 35 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x37
timestamp 1713382353
transform 1 0 36 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x38
timestamp 1713382353
transform 1 0 37 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x39
timestamp 1713382353
transform 1 0 38 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x40
timestamp 1713382353
transform 1 0 39 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x41
timestamp 1713382353
transform 1 0 40 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x42
timestamp 1713382353
transform 1 0 41 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x43
timestamp 1713382353
transform 1 0 42 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x44
timestamp 1713382353
transform 1 0 43 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x45
timestamp 1713382353
transform 1 0 44 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x46
timestamp 1713382353
transform 1 0 45 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x47
timestamp 1713382353
transform 1 0 46 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x48
timestamp 1713382353
transform 1 0 47 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x49
timestamp 1713382353
transform 1 0 48 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x50
timestamp 1713382353
transform 1 0 49 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x51
timestamp 1713382353
transform 1 0 50 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x52
timestamp 1713382353
transform 1 0 51 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x53
timestamp 1713382353
transform 1 0 52 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x54
timestamp 1713382353
transform 1 0 53 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x55
timestamp 1713382353
transform 1 0 54 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x56
timestamp 1713382353
transform 1 0 55 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x57
timestamp 1713382353
transform 1 0 56 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x58
timestamp 1713382353
transform 1 0 57 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x59
timestamp 1713382353
transform 1 0 58 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x60
timestamp 1713382353
transform 1 0 59 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x61
timestamp 1713382353
transform 1 0 60 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x62
timestamp 1713382353
transform 1 0 61 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x63
timestamp 1713382353
transform 1 0 62 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x64
timestamp 1713382353
transform 1 0 63 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x65
timestamp 1713382353
transform 1 0 64 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x66
timestamp 1713382353
transform 1 0 65 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x67
timestamp 1713382353
transform 1 0 66 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x68
timestamp 1713382353
transform 1 0 67 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x69
timestamp 1713382353
transform 1 0 68 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x70
timestamp 1713382353
transform 1 0 69 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x71
timestamp 1713382353
transform 1 0 70 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x72
timestamp 1713382353
transform 1 0 71 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x73
timestamp 1713382353
transform 1 0 72 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x74
timestamp 1713382353
transform 1 0 73 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x75
timestamp 1713382353
transform 1 0 74 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x76
timestamp 1713382353
transform 1 0 75 0 1 600
box -53 -1200 611 3001
use SUNTR_NCHLCM  x77
timestamp 1713382353
transform 1 0 76 0 1 600
box -53 -1200 1611 2983
use SUNTR_PCHLCM  x78
timestamp 1713382353
transform 1 0 77 0 1 600
box -53 -1200 611 3001
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD_1V8
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Clk
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Clk_1
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Clk_2
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
