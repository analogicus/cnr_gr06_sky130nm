*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR06_main_lpe.spi
#else
.include ../../../work/xsch/CNR_GR06_main.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS (Common for all corners)
*-----------------------------------------------------------------
.param TRF = 100p
.param t_start = 0.5u
.param t_start_del = {t_start + TRF}
.param PERIOD_CLK = 500n
.param PW_CLK = PERIOD_CLK/2
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0  dc 0
VDD  VDD_1V8 0 dc 1.2
Vdref Vdref 0 dc 1.2
VT2  VT2 0 SIN(0 0.25 10000 0 0 180)
VT1  VT1 0 SIN(0 0.25 10000 0 0)
VBP VBP 0 dc 0.08
VBN VBN 0 dc 1.12
VCLK Clk 0 dc 0 pulse 0 1.2 {t_start} {TRF} {TRF} {PW_CLK} {PERIOD_CLK}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*-----------------------------------------------------------------
* PROBE
*-----------------------------------------------------------------
#ifdef Debug
.save all
#else
.save ${VPORTS}
#endif

*-----------------------------------------------------------------
* NGSPICE control - Corner Simulation Example
*-----------------------------------------------------------------
.control
* Run the simulation for fast corner
set param vth0_n=0.47
set param vth0_p=-0.47
run
set filetype=ascii
write output_data_fast.txt V(Voc)

* Run the simulation for slow corner
set param vth0_n=0.53
set param vth0_p=-0.53
run
set filetype=ascii
write output_data_slow.txt V(Voc)
.endc

.end

