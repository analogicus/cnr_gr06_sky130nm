*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR06_lpe.spi
#else
.include ../../../work/xsch/CNR_GR06.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

.param TRF = 100p

.param t_start = 0.5u
.param t_start_del = {t_start + TRF}

*- 8 MHz clock frequency
.param PERIOD_CLK = 0.5u

*- 25% duty-cycle clock
.param PW_CLK = PERIOD_CLK/2
*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0  dc 0
VDD  VDD_1V8 0 dc {AVDD}
Vref Vref 0 dc 0.2

VCLK Clk 0 dc 0 pulse 0 1.8 {t_start} {TRF} {TRF} {PW_CLK} {PERIOD_CLK}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save ${VPORTS}
#endif

*.save v(vp,vn)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 10n 10u 0

tran 1n 10u
write
quit

.endc

.end
