*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR06_main_lpe.spi
#else
.include ../../../work/xsch/CNR_GR06_main.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 100p

.param t_start = 0.5u
.param t_start_del = {t_start + TRF}

*- 8 MHz clock frequency
*.param PERIOD_CLK = 250n

*- 25% duty-cycle clock
*.param PW_CLK = PERIOD_CLK/2

*- Supply, vdda is set in includes
.param AVDD = {vdda}
*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0  dc 0
VDD  VDD_1V8 0 dc {AVDD}
Vdref Vdref 0 dc 0.8

*VT2 VT2 0 dc 0.2
*VT1 VT1 0 dc 1.2

VT2  VT2 0 SIN(0.6 0.6 50000 0 0 180)
VT1  VT1 0 SIN(0.6 0.6 50000 0 0)

*VCLK Clk 0 dc 0 pulse 0 {AVDD} {t_start} {TRF} {TRF} {PW_CLK} {PERIOD_CLK}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save ${VPORTS}
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 1 1 1 10n 1u 0

dc TEMP -40 125 5
write
quit

.endc

.end
