magic
tech sky130B
magscale 1 2
timestamp 1713381639
<< checkpaint >>
rect -1260 -8060 1460 1460
rect 1679 -1361977 11450 -1361177
rect -1260 -1368864 14389 -1361977
<< error_p >>
rect 20629 1204800 20630 1210881
rect 27001 945560 27002 951641
rect 33373 781120 33374 787201
rect 39745 521920 39746 527961
rect 46117 262640 46118 268721
rect 54318 11009 54353 11043
rect 54319 10990 54353 11009
rect 54338 10735 54353 10990
rect 54372 10956 54407 10990
rect 54857 10956 54892 10990
rect 54372 10735 54406 10956
rect 54858 10937 54892 10956
rect 54877 10735 54892 10937
rect 54911 10903 54946 10937
rect 55396 10903 55431 10937
rect 54911 10735 54945 10903
rect 55397 10884 55431 10903
rect 55416 10735 55431 10884
rect 55450 10850 55485 10884
rect 55935 10850 55970 10884
rect 55450 10735 55484 10850
rect 55936 10831 55970 10850
rect 55955 10735 55970 10831
rect 55989 10797 56024 10831
rect 55989 10735 56023 10797
rect 52668 6800 52690 7000
rect 52696 6800 52718 7000
rect 52869 6800 52896 7000
rect 52897 6800 52924 7000
rect 53070 6800 53097 7000
rect 53098 6800 53125 7000
rect 53271 6800 53298 7000
rect 53299 6800 53326 7000
rect 53477 6800 53499 7000
rect 53505 6800 53527 7000
rect 53683 6800 53705 7000
rect 53711 6800 53733 7000
rect 53884 6800 53911 7000
rect 53912 6800 53939 7000
rect 54085 6800 54112 7000
rect 54113 6800 54140 7000
rect 54291 6800 54313 7000
rect 54319 6800 54341 7000
rect 54497 6800 54519 7000
rect 54525 6800 54547 7000
rect 54703 6800 54725 7000
rect 54731 6800 54753 7000
rect 54904 6800 54931 7000
rect 54932 6800 54959 7000
rect 55110 6800 55132 7000
rect 55138 6800 55160 7000
rect 55311 6800 55338 7000
rect 55339 6800 55366 7000
rect 55517 6800 55539 7000
rect 55545 6800 55567 7000
rect 55718 6800 55745 7000
rect 55746 6800 55773 7000
rect 55924 6800 55946 7000
rect 55952 6800 55974 7000
rect 56125 6800 56152 7000
rect 56153 6800 56180 7000
rect 56331 6800 56353 7000
rect 56359 6800 56381 7000
rect 56532 6800 56559 7000
rect 56560 6800 56587 7000
rect 56738 6800 56760 7000
rect 56766 6800 56788 7000
rect 56944 6800 56966 7000
rect 56972 6800 56994 7000
rect 57145 6800 57172 7000
rect 57173 6800 57200 7000
rect 57346 6800 57373 7000
rect 57374 6800 57401 7000
rect 57552 6800 57574 7000
rect 57580 6800 57602 7000
rect 57753 6800 57780 7000
rect 57781 6800 57808 7000
rect 57959 6800 57981 7000
rect 57987 6800 58009 7000
rect 58160 6800 58187 7000
rect 58188 6800 58215 7000
rect 58366 6800 58388 7000
rect 58394 6800 58416 7000
rect 58567 6800 58594 7000
rect 58595 6800 58622 7000
rect 58773 6800 58795 7000
rect 58801 6800 58823 7000
rect 58974 6800 59001 7000
rect 59002 6800 59029 7000
rect 59180 6800 59202 7000
rect 59208 6800 59230 7000
rect 59381 6800 59408 7000
rect 59409 6800 59436 7000
rect 59587 6800 59609 7000
rect 59615 6800 59637 7000
rect 59788 6800 59815 7000
rect 59816 6800 59843 7000
rect 59994 6800 60016 7000
rect 60022 6800 60044 7000
rect 60195 6800 60222 7000
rect 60223 6800 60250 7000
rect 60401 6800 60423 7000
rect 60429 6800 60451 7000
rect 72556 6903 72591 6937
rect 72557 6884 72591 6903
rect 52668 6400 52690 6600
rect 52696 6400 52718 6600
rect 52869 6400 52896 6600
rect 52897 6400 52924 6600
rect 53070 6400 53097 6600
rect 53098 6400 53125 6600
rect 53271 6400 53298 6600
rect 53299 6400 53326 6600
rect 53477 6400 53499 6600
rect 53505 6400 53527 6600
rect 53683 6400 53705 6600
rect 53711 6400 53733 6600
rect 53884 6400 53911 6600
rect 53912 6400 53939 6600
rect 54085 6400 54112 6600
rect 54113 6400 54140 6600
rect 54291 6400 54313 6600
rect 54319 6400 54341 6600
rect 54497 6400 54519 6600
rect 54525 6400 54547 6600
rect 54703 6400 54725 6600
rect 54731 6400 54753 6600
rect 54904 6400 54931 6600
rect 54932 6400 54959 6600
rect 55110 6400 55132 6600
rect 55138 6400 55160 6600
rect 55311 6400 55338 6600
rect 55339 6400 55366 6600
rect 55517 6400 55539 6600
rect 55545 6400 55567 6600
rect 55718 6400 55745 6600
rect 55746 6400 55773 6600
rect 55924 6400 55946 6600
rect 55952 6400 55974 6600
rect 56125 6400 56152 6600
rect 56153 6400 56180 6600
rect 56331 6400 56353 6600
rect 56359 6400 56381 6600
rect 56532 6400 56559 6600
rect 56560 6400 56587 6600
rect 56738 6400 56760 6600
rect 56766 6400 56788 6600
rect 56944 6400 56966 6600
rect 56972 6400 56994 6600
rect 57145 6400 57172 6600
rect 57173 6400 57200 6600
rect 57346 6400 57373 6600
rect 57374 6400 57401 6600
rect 57552 6400 57574 6600
rect 57580 6400 57602 6600
rect 57753 6400 57780 6600
rect 57781 6400 57808 6600
rect 57959 6400 57981 6600
rect 57987 6400 58009 6600
rect 58160 6400 58187 6600
rect 58188 6400 58215 6600
rect 58366 6400 58388 6600
rect 58394 6400 58416 6600
rect 58567 6400 58594 6600
rect 58595 6400 58622 6600
rect 58773 6400 58795 6600
rect 58801 6400 58823 6600
rect 58974 6400 59001 6600
rect 59002 6400 59029 6600
rect 59180 6400 59202 6600
rect 59208 6400 59230 6600
rect 59381 6400 59408 6600
rect 59409 6400 59436 6600
rect 59587 6400 59609 6600
rect 59615 6400 59637 6600
rect 59788 6400 59815 6600
rect 59816 6400 59843 6600
rect 59994 6400 60016 6600
rect 60022 6400 60044 6600
rect 60195 6400 60222 6600
rect 60223 6400 60250 6600
rect 60401 6400 60423 6600
rect 60429 6400 60451 6600
rect 71478 4991 71513 5025
rect 72071 5008 72105 5026
rect 71479 4972 71513 4991
rect 71498 2677 71513 4972
rect 71532 4938 71567 4972
rect 71532 2677 71566 4938
rect 71532 2643 71547 2677
rect 72035 2624 72105 5008
rect 72035 2588 72088 2624
rect 72576 2571 72591 6884
rect 72610 6850 72645 6884
rect 72610 2571 72644 6850
rect 72610 2537 72625 2571
rect 21977 997 22012 1031
rect 21978 978 22012 997
rect 21997 583 22012 978
rect 22031 944 22066 978
rect 22516 944 22551 978
rect 22031 583 22065 944
rect 22517 925 22551 944
rect 22031 549 22046 583
rect 22536 530 22551 925
rect 22570 891 22605 925
rect 23055 891 23090 925
rect 22570 530 22604 891
rect 23056 872 23090 891
rect 22570 496 22585 530
rect 23075 477 23090 872
rect 23109 838 23144 872
rect 23594 838 23629 872
rect 23109 477 23143 838
rect 23595 819 23629 838
rect 23109 443 23124 477
rect 23614 424 23629 819
rect 23648 785 23683 819
rect 24133 785 24168 819
rect 23648 424 23682 785
rect 24134 766 24168 785
rect 23648 390 23663 424
rect 24153 371 24168 766
rect 24187 732 24222 766
rect 24672 732 24707 766
rect 24187 371 24221 732
rect 24673 713 24707 732
rect 24187 337 24202 371
rect 24692 318 24707 713
rect 24726 679 24761 713
rect 24726 318 24760 679
rect 24726 284 24741 318
rect 6371 -163240 6373 -157159
rect 12743 -422480 12745 -416399
rect 19115 -586920 19117 -580839
rect 25487 -846120 25489 -840079
rect 31859 -1105400 31861 -1099319
rect 59583 -1360231 59618 -1360197
rect 59584 -1360250 59618 -1360231
rect 59603 -1364563 59618 -1360250
rect 59637 -1360284 59672 -1360250
rect 60122 -1360284 60157 -1360250
rect 59637 -1364563 59671 -1360284
rect 60123 -1360303 60157 -1360284
rect 59637 -1364597 59652 -1364563
rect 60142 -1364616 60157 -1360303
rect 60176 -1360337 60211 -1360303
rect 60661 -1360337 60696 -1360303
rect 60176 -1364616 60210 -1360337
rect 60662 -1360356 60696 -1360337
rect 60176 -1364650 60191 -1364616
rect 60681 -1364669 60696 -1360356
rect 60715 -1360390 60750 -1360356
rect 61200 -1360390 61235 -1360356
rect 60715 -1364669 60749 -1360390
rect 61201 -1360409 61235 -1360390
rect 60715 -1364703 60730 -1364669
rect 61220 -1364722 61235 -1360409
rect 61254 -1360443 61289 -1360409
rect 61739 -1360443 61774 -1360409
rect 61254 -1364722 61288 -1360443
rect 61740 -1360462 61774 -1360443
rect 61254 -1364756 61269 -1364722
rect 61759 -1364775 61774 -1360462
rect 61793 -1360496 61828 -1360462
rect 61793 -1364775 61827 -1360496
rect 67912 -1361137 67947 -1361103
rect 67913 -1361156 67947 -1361137
rect 62279 -1362497 62313 -1362479
rect 62279 -1362533 62349 -1362497
rect 62296 -1362567 62367 -1362533
rect 62817 -1362567 62852 -1362533
rect 61793 -1364809 61808 -1364775
rect 62296 -1364828 62366 -1362567
rect 62818 -1362586 62852 -1362567
rect 62296 -1364864 62349 -1364828
rect 62837 -1364881 62852 -1362586
rect 62871 -1362620 62906 -1362586
rect 63356 -1362620 63391 -1362586
rect 63949 -1362603 63983 -1362585
rect 62871 -1364881 62905 -1362620
rect 63357 -1362639 63391 -1362620
rect 62871 -1364915 62886 -1364881
rect 63376 -1364934 63391 -1362639
rect 63410 -1362673 63445 -1362639
rect 63410 -1364934 63444 -1362673
rect 63410 -1364968 63425 -1364934
rect 63913 -1364987 63983 -1362603
rect 64435 -1362709 64469 -1362691
rect 64435 -1362745 64505 -1362709
rect 64452 -1362779 64523 -1362745
rect 64973 -1362779 65008 -1362745
rect 63913 -1365023 63966 -1364987
rect 64452 -1365040 64522 -1362779
rect 64974 -1362798 65008 -1362779
rect 64452 -1365076 64505 -1365040
rect 64993 -1365093 65008 -1362798
rect 65027 -1362832 65062 -1362798
rect 65027 -1365093 65061 -1362832
rect 65757 -1362926 65791 -1362908
rect 65757 -1362962 65827 -1362926
rect 65774 -1362996 65845 -1362962
rect 66295 -1362996 66330 -1362962
rect 65027 -1365127 65042 -1365093
rect 65774 -1365257 65844 -1362996
rect 66296 -1363015 66330 -1362996
rect 65774 -1365293 65827 -1365257
rect 66315 -1365310 66330 -1363015
rect 66349 -1363049 66384 -1363015
rect 66834 -1363049 66869 -1363015
rect 67427 -1363032 67461 -1363014
rect 66349 -1365310 66383 -1363049
rect 66835 -1363068 66869 -1363049
rect 66349 -1365344 66364 -1365310
rect 66854 -1365363 66869 -1363068
rect 66888 -1363102 66923 -1363068
rect 66888 -1365363 66922 -1363102
rect 66888 -1365397 66903 -1365363
rect 67391 -1365416 67461 -1363032
rect 67391 -1365452 67444 -1365416
rect 67932 -1365469 67947 -1361156
rect 67966 -1361190 68001 -1361156
rect 67966 -1365469 68000 -1361190
rect 67966 -1365503 67981 -1365469
<< error_s >>
rect 60602 6800 60629 7000
rect 60630 6800 60657 7000
rect 60808 6800 60830 7000
rect 60836 6800 60858 7000
rect 61009 6800 61036 7000
rect 61037 6800 61064 7000
rect 61215 6800 61237 7000
rect 61243 6800 61265 7000
rect 61416 6800 61443 7000
rect 61444 6800 61471 7000
rect 61622 6800 61644 7000
rect 61650 6800 61672 7000
rect 61823 6800 61850 7000
rect 61851 6800 61878 7000
rect 62029 6800 62051 7000
rect 62057 6800 62079 7000
rect 62230 6800 62257 7000
rect 62258 6800 62285 7000
rect 62436 6800 62458 7000
rect 62464 6800 62486 7000
rect 62637 6800 62664 7000
rect 62665 6800 62692 7000
rect 62843 6800 62865 7000
rect 62871 6800 62893 7000
rect 63044 6800 63071 7000
rect 63072 6800 63099 7000
rect 63250 6800 63272 7000
rect 63278 6800 63300 7000
rect 63451 6800 63478 7000
rect 63479 6800 63506 7000
rect 63657 6800 63679 7000
rect 63685 6800 63707 7000
rect 63858 6800 63885 7000
rect 63886 6800 63913 7000
rect 64064 6800 64086 7000
rect 64092 6800 64114 7000
rect 64265 6800 64292 7000
rect 64293 6800 64320 7000
rect 64471 6800 64493 7000
rect 64499 6800 64521 7000
rect 64672 6800 64699 7000
rect 64700 6800 64727 7000
rect 64878 6800 64900 7000
rect 64906 6800 64928 7000
rect 65079 6800 65106 7000
rect 65107 6800 65134 7000
rect 65285 6800 65307 7000
rect 65313 6800 65335 7000
rect 65486 6800 65513 7000
rect 65514 6800 65541 7000
rect 65692 6800 65714 7000
rect 65720 6800 65742 7000
rect 65893 6800 65920 7000
rect 65921 6800 65948 7000
rect 66099 6800 66121 7000
rect 66127 6800 66149 7000
rect 66300 6800 66327 7000
rect 66328 6800 66355 7000
rect 66506 6800 66528 7000
rect 66534 6800 66556 7000
rect 66707 6800 66734 7000
rect 66735 6800 66762 7000
rect 66913 6800 66935 7000
rect 66941 6800 66963 7000
rect 67114 6800 67141 7000
rect 67142 6800 67169 7000
rect 67320 6800 67342 7000
rect 67348 6800 67370 7000
rect 67521 6800 67548 7000
rect 67549 6800 67576 7000
rect 67727 6800 67749 7000
rect 67755 6800 67777 7000
rect 67928 6800 67955 7000
rect 67956 6800 67983 7000
rect 68134 6800 68156 7000
rect 68162 6800 68184 7000
rect 60602 6400 60629 6600
rect 60630 6400 60657 6600
rect 60808 6400 60830 6600
rect 60836 6400 60858 6600
rect 61009 6400 61036 6600
rect 61037 6400 61064 6600
rect 61215 6400 61237 6600
rect 61243 6400 61265 6600
rect 61416 6400 61443 6600
rect 61444 6400 61471 6600
rect 61622 6400 61644 6600
rect 61650 6400 61672 6600
rect 61823 6400 61850 6600
rect 61851 6400 61878 6600
rect 62029 6400 62051 6600
rect 62057 6400 62079 6600
rect 62230 6400 62257 6600
rect 62258 6400 62285 6600
rect 62436 6400 62458 6600
rect 62464 6400 62486 6600
rect 62637 6400 62664 6600
rect 62665 6400 62692 6600
rect 62843 6400 62865 6600
rect 62871 6400 62893 6600
rect 63044 6400 63071 6600
rect 63072 6400 63099 6600
rect 63250 6400 63272 6600
rect 63278 6400 63300 6600
rect 63451 6400 63478 6600
rect 63479 6400 63506 6600
rect 63657 6400 63679 6600
rect 63685 6400 63707 6600
rect 63858 6400 63885 6600
rect 63886 6400 63913 6600
rect 64064 6400 64086 6600
rect 64092 6400 64114 6600
rect 64265 6400 64292 6600
rect 64293 6400 64320 6600
rect 64471 6400 64493 6600
rect 64499 6400 64521 6600
rect 64672 6400 64699 6600
rect 64700 6400 64727 6600
rect 64878 6400 64900 6600
rect 64906 6400 64928 6600
rect 65079 6400 65106 6600
rect 65107 6400 65134 6600
rect 65285 6400 65307 6600
rect 65313 6400 65335 6600
rect 65486 6400 65513 6600
rect 65514 6400 65541 6600
rect 65692 6400 65714 6600
rect 65720 6400 65742 6600
rect 65893 6400 65920 6600
rect 65921 6400 65948 6600
rect 66099 6400 66121 6600
rect 66127 6400 66149 6600
rect 66300 6400 66327 6600
rect 66328 6400 66355 6600
rect 66506 6400 66528 6600
rect 66534 6400 66556 6600
rect 66707 6400 66734 6600
rect 66735 6400 66762 6600
rect 66913 6400 66935 6600
rect 66941 6400 66963 6600
rect 67114 6400 67141 6600
rect 67142 6400 67169 6600
rect 67320 6400 67342 6600
rect 67348 6400 67370 6600
rect 67521 6400 67548 6600
rect 67549 6400 67576 6600
rect 67727 6400 67749 6600
rect 67755 6400 67777 6600
rect 67928 6400 67955 6600
rect 67956 6400 67983 6600
rect 68134 6400 68156 6600
rect 68162 6400 68184 6600
rect 52668 6000 52690 6200
rect 52696 6000 52718 6200
rect 52869 6000 52896 6200
rect 52897 6000 52924 6200
rect 53070 6000 53097 6200
rect 53098 6000 53125 6200
rect 53271 6000 53298 6200
rect 53299 6000 53326 6200
rect 53477 6000 53499 6200
rect 53505 6000 53527 6200
rect 53683 6000 53705 6200
rect 53711 6000 53733 6200
rect 53884 6000 53911 6200
rect 53912 6000 53939 6200
rect 54085 6000 54112 6200
rect 54113 6000 54140 6200
rect 54291 6000 54313 6200
rect 54319 6000 54341 6200
rect 54497 6000 54519 6200
rect 54525 6000 54547 6200
rect 54703 6000 54725 6200
rect 54731 6000 54753 6200
rect 54904 6000 54931 6200
rect 54932 6000 54959 6200
rect 55110 6000 55132 6200
rect 55138 6000 55160 6200
rect 55311 6000 55338 6200
rect 55339 6000 55366 6200
rect 55517 6000 55539 6200
rect 55545 6000 55567 6200
rect 55718 6000 55745 6200
rect 55746 6000 55773 6200
rect 55924 6000 55946 6200
rect 55952 6000 55974 6200
rect 56125 6000 56152 6200
rect 56153 6000 56180 6200
rect 56331 6000 56353 6200
rect 56359 6000 56381 6200
rect 56532 6000 56559 6200
rect 56560 6000 56587 6200
rect 56738 6000 56760 6200
rect 56766 6000 56788 6200
rect 56944 6000 56966 6200
rect 56972 6000 56994 6200
rect 57145 6000 57172 6200
rect 57173 6000 57200 6200
rect 57346 6000 57373 6200
rect 57374 6000 57401 6200
rect 57552 6000 57574 6200
rect 57580 6000 57602 6200
rect 57753 6000 57780 6200
rect 57781 6000 57808 6200
rect 57959 6000 57981 6200
rect 57987 6000 58009 6200
rect 58160 6000 58187 6200
rect 58188 6000 58215 6200
rect 58366 6000 58388 6200
rect 58394 6000 58416 6200
rect 58567 6000 58594 6200
rect 58595 6000 58622 6200
rect 58773 6000 58795 6200
rect 58801 6000 58823 6200
rect 58974 6000 59001 6200
rect 59002 6000 59029 6200
rect 59180 6000 59202 6200
rect 59208 6000 59230 6200
rect 59381 6000 59408 6200
rect 59409 6000 59436 6200
rect 59587 6000 59609 6200
rect 59615 6000 59637 6200
rect 59788 6000 59815 6200
rect 59816 6000 59843 6200
rect 59994 6000 60016 6200
rect 60022 6000 60044 6200
rect 60195 6000 60222 6200
rect 60223 6000 60250 6200
rect 60401 6000 60423 6200
rect 60429 6000 60451 6200
rect 60602 6000 60629 6200
rect 60630 6000 60657 6200
rect 60808 6000 60830 6200
rect 60836 6000 60858 6200
rect 61009 6000 61036 6200
rect 61037 6000 61064 6200
rect 61215 6000 61237 6200
rect 61243 6000 61265 6200
rect 61416 6000 61443 6200
rect 61444 6000 61471 6200
rect 61622 6000 61644 6200
rect 61650 6000 61672 6200
rect 61823 6000 61850 6200
rect 61851 6000 61878 6200
rect 62029 6000 62051 6200
rect 62057 6000 62079 6200
rect 62230 6000 62257 6200
rect 62258 6000 62285 6200
rect 62436 6000 62458 6200
rect 62464 6000 62486 6200
rect 62637 6000 62664 6200
rect 62665 6000 62692 6200
rect 62843 6000 62865 6200
rect 62871 6000 62893 6200
rect 63044 6000 63071 6200
rect 63072 6000 63099 6200
rect 63250 6000 63272 6200
rect 63278 6000 63300 6200
rect 63451 6000 63478 6200
rect 63479 6000 63506 6200
rect 63657 6000 63679 6200
rect 63685 6000 63707 6200
rect 63858 6000 63885 6200
rect 63886 6000 63913 6200
rect 64064 6000 64086 6200
rect 64092 6000 64114 6200
rect 64265 6000 64292 6200
rect 64293 6000 64320 6200
rect 64471 6000 64493 6200
rect 64499 6000 64521 6200
rect 64672 6000 64699 6200
rect 64700 6000 64727 6200
rect 64878 6000 64900 6200
rect 64906 6000 64928 6200
rect 65079 6000 65106 6200
rect 65107 6000 65134 6200
rect 65285 6000 65307 6200
rect 65313 6000 65335 6200
rect 65486 6000 65513 6200
rect 65514 6000 65541 6200
rect 65692 6000 65714 6200
rect 65720 6000 65742 6200
rect 65893 6000 65920 6200
rect 65921 6000 65948 6200
rect 66099 6000 66121 6200
rect 66127 6000 66149 6200
rect 66300 6000 66327 6200
rect 66328 6000 66355 6200
rect 66506 6000 66528 6200
rect 66534 6000 66556 6200
rect 66707 6000 66734 6200
rect 66735 6000 66762 6200
rect 66913 6000 66935 6200
rect 66941 6000 66963 6200
rect 67114 6000 67141 6200
rect 67142 6000 67169 6200
rect 67320 6000 67342 6200
rect 67348 6000 67370 6200
rect 67521 6000 67548 6200
rect 67549 6000 67576 6200
rect 67727 6000 67749 6200
rect 67755 6000 67777 6200
rect 67928 6000 67955 6200
rect 67956 6000 67983 6200
rect 68134 6000 68156 6200
rect 68162 6000 68184 6200
rect 52869 5600 52896 5800
rect 52897 5600 52924 5800
rect 53070 5600 53097 5800
rect 53098 5600 53125 5800
rect 53271 5600 53298 5800
rect 53299 5600 53326 5800
rect 53477 5600 53499 5800
rect 53505 5600 53527 5800
rect 53683 5600 53705 5800
rect 53711 5600 53733 5800
rect 53884 5600 53911 5800
rect 53912 5600 53939 5800
rect 54085 5600 54112 5800
rect 54113 5600 54140 5800
rect 54291 5600 54313 5800
rect 54319 5600 54341 5800
rect 54497 5600 54519 5800
rect 54525 5600 54547 5800
rect 54703 5600 54725 5800
rect 54731 5600 54753 5800
rect 54904 5600 54931 5800
rect 54932 5600 54959 5800
rect 55110 5600 55132 5800
rect 55138 5600 55160 5800
rect 55311 5600 55338 5800
rect 55339 5600 55366 5800
rect 55517 5600 55539 5800
rect 55545 5600 55567 5800
rect 55718 5600 55745 5800
rect 55746 5600 55773 5800
rect 55924 5600 55946 5800
rect 55952 5600 55974 5800
rect 56125 5600 56152 5800
rect 56153 5600 56180 5800
rect 56331 5600 56353 5800
rect 56359 5600 56381 5800
rect 56532 5600 56559 5800
rect 56560 5600 56587 5800
rect 56738 5600 56760 5800
rect 56766 5600 56788 5800
rect 56944 5600 56966 5800
rect 56972 5600 56994 5800
rect 57145 5600 57172 5800
rect 57173 5600 57200 5800
rect 57346 5600 57373 5800
rect 57374 5600 57401 5800
rect 57552 5600 57574 5800
rect 57580 5600 57602 5800
rect 57753 5600 57780 5800
rect 57781 5600 57808 5800
rect 57959 5600 57981 5800
rect 57987 5600 58009 5800
rect 58160 5600 58187 5800
rect 58188 5600 58215 5800
rect 58366 5600 58388 5800
rect 58394 5600 58416 5800
rect 58567 5600 58594 5800
rect 58595 5600 58622 5800
rect 58773 5600 58795 5800
rect 58801 5600 58823 5800
rect 58974 5600 59001 5800
rect 59002 5600 59029 5800
rect 59180 5600 59202 5800
rect 59208 5600 59230 5800
rect 59381 5600 59408 5800
rect 59409 5600 59436 5800
rect 59587 5600 59609 5800
rect 59615 5600 59637 5800
rect 59788 5600 59815 5800
rect 59816 5600 59843 5800
rect 59994 5600 60016 5800
rect 60022 5600 60044 5800
rect 60195 5600 60222 5800
rect 60223 5600 60250 5800
rect 60401 5600 60423 5800
rect 60429 5600 60451 5800
rect 60602 5600 60629 5800
rect 60630 5600 60657 5800
rect 60808 5600 60830 5800
rect 60836 5600 60858 5800
rect 61009 5600 61036 5800
rect 61037 5600 61064 5800
rect 61215 5600 61237 5800
rect 61243 5600 61265 5800
rect 61416 5600 61443 5800
rect 61444 5600 61471 5800
rect 61622 5600 61644 5800
rect 61650 5600 61672 5800
rect 61823 5600 61850 5800
rect 61851 5600 61878 5800
rect 62029 5600 62051 5800
rect 62057 5600 62079 5800
rect 62230 5600 62257 5800
rect 62258 5600 62285 5800
rect 62436 5600 62458 5800
rect 62464 5600 62486 5800
rect 62637 5600 62664 5800
rect 62665 5600 62692 5800
rect 62843 5600 62865 5800
rect 62871 5600 62893 5800
rect 63044 5600 63071 5800
rect 63072 5600 63099 5800
rect 63250 5600 63272 5800
rect 63278 5600 63300 5800
rect 63451 5600 63478 5800
rect 63479 5600 63506 5800
rect 63657 5600 63679 5800
rect 63685 5600 63707 5800
rect 63858 5600 63885 5800
rect 63886 5600 63913 5800
rect 64064 5600 64086 5800
rect 64092 5600 64114 5800
rect 64265 5600 64292 5800
rect 64293 5600 64320 5800
rect 64471 5600 64493 5800
rect 64499 5600 64521 5800
rect 64672 5600 64699 5800
rect 64700 5600 64727 5800
rect 64878 5600 64900 5800
rect 64906 5600 64928 5800
rect 65079 5600 65106 5800
rect 65107 5600 65134 5800
rect 65285 5600 65307 5800
rect 65313 5600 65335 5800
rect 65486 5600 65513 5800
rect 65514 5600 65541 5800
rect 65692 5600 65714 5800
rect 65720 5600 65742 5800
rect 65893 5600 65920 5800
rect 65921 5600 65948 5800
rect 66099 5600 66121 5800
rect 66127 5600 66149 5800
rect 66300 5600 66327 5800
rect 66328 5600 66355 5800
rect 66506 5600 66528 5800
rect 66534 5600 66556 5800
rect 66707 5600 66734 5800
rect 66735 5600 66762 5800
rect 66913 5600 66935 5800
rect 66941 5600 66963 5800
rect 67114 5600 67141 5800
rect 67142 5600 67169 5800
rect 67320 5600 67342 5800
rect 67348 5600 67370 5800
rect 67521 5600 67548 5800
rect 67549 5600 67576 5800
rect 67727 5600 67749 5800
rect 67755 5600 67777 5800
rect 67928 5600 67955 5800
rect 67956 5600 67983 5800
rect 68134 5600 68156 5800
rect 68162 5600 68184 5800
rect 52869 5200 52896 5400
rect 52897 5200 52924 5400
rect 53070 5200 53097 5400
rect 53098 5200 53125 5400
rect 53271 5200 53298 5400
rect 53299 5200 53326 5400
rect 53477 5200 53499 5400
rect 53505 5200 53527 5400
rect 53683 5200 53705 5400
rect 53711 5200 53733 5400
rect 53884 5200 53911 5400
rect 53912 5200 53939 5400
rect 54085 5200 54112 5400
rect 54113 5200 54140 5400
rect 54291 5200 54313 5400
rect 54319 5200 54341 5400
rect 54497 5200 54519 5400
rect 54525 5200 54547 5400
rect 54703 5200 54725 5400
rect 54731 5200 54753 5400
rect 54904 5200 54931 5400
rect 54932 5200 54959 5400
rect 55110 5200 55132 5400
rect 55138 5200 55160 5400
rect 55311 5200 55338 5400
rect 55339 5200 55366 5400
rect 55517 5200 55539 5400
rect 55545 5200 55567 5400
rect 55718 5200 55745 5400
rect 55746 5200 55773 5400
rect 55924 5200 55946 5400
rect 55952 5200 55974 5400
rect 56125 5200 56152 5400
rect 56153 5200 56180 5400
rect 56331 5200 56353 5400
rect 56359 5200 56381 5400
rect 56532 5200 56559 5400
rect 56560 5200 56587 5400
rect 56738 5200 56760 5400
rect 56766 5200 56788 5400
rect 56944 5200 56966 5400
rect 56972 5200 56994 5400
rect 57145 5200 57172 5400
rect 57173 5200 57200 5400
rect 57346 5200 57373 5400
rect 57374 5200 57401 5400
rect 57552 5200 57574 5400
rect 57580 5200 57602 5400
rect 57753 5200 57780 5400
rect 57781 5200 57808 5400
rect 57959 5200 57981 5400
rect 57987 5200 58009 5400
rect 58160 5200 58187 5400
rect 58188 5200 58215 5400
rect 58366 5200 58388 5400
rect 58394 5200 58416 5400
rect 58567 5200 58594 5400
rect 58595 5200 58622 5400
rect 58773 5200 58795 5400
rect 58801 5200 58823 5400
rect 58974 5200 59001 5400
rect 59002 5200 59029 5400
rect 59180 5200 59202 5400
rect 59208 5200 59230 5400
rect 59381 5200 59408 5400
rect 59409 5200 59436 5400
rect 59587 5200 59609 5400
rect 59615 5200 59637 5400
rect 59788 5200 59815 5400
rect 59816 5200 59843 5400
rect 59994 5200 60016 5400
rect 60022 5200 60044 5400
rect 60195 5200 60222 5400
rect 60223 5200 60250 5400
rect 60401 5200 60423 5400
rect 60429 5200 60451 5400
rect 60602 5200 60629 5400
rect 60630 5200 60657 5400
rect 60808 5200 60830 5400
rect 60836 5200 60858 5400
rect 61009 5200 61036 5400
rect 61037 5200 61064 5400
rect 61215 5200 61237 5400
rect 61243 5200 61265 5400
rect 61416 5200 61443 5400
rect 61444 5200 61471 5400
rect 61622 5200 61644 5400
rect 61650 5200 61672 5400
rect 61823 5200 61850 5400
rect 61851 5200 61878 5400
rect 62029 5200 62051 5400
rect 62057 5200 62079 5400
rect 62230 5200 62257 5400
rect 62258 5200 62285 5400
rect 62436 5200 62458 5400
rect 62464 5200 62486 5400
rect 62637 5200 62664 5400
rect 62665 5200 62692 5400
rect 62843 5200 62865 5400
rect 62871 5200 62893 5400
rect 63044 5200 63071 5400
rect 63072 5200 63099 5400
rect 63250 5200 63272 5400
rect 63278 5200 63300 5400
rect 63451 5200 63478 5400
rect 63479 5200 63506 5400
rect 63657 5200 63679 5400
rect 63685 5200 63707 5400
rect 63858 5200 63885 5400
rect 63886 5200 63913 5400
rect 64064 5200 64086 5400
rect 64092 5200 64114 5400
rect 64265 5200 64292 5400
rect 64293 5200 64320 5400
rect 64471 5200 64493 5400
rect 64499 5200 64521 5400
rect 64672 5200 64699 5400
rect 64700 5200 64727 5400
rect 64878 5200 64900 5400
rect 64906 5200 64928 5400
rect 65079 5200 65106 5400
rect 65107 5200 65134 5400
rect 65285 5200 65307 5400
rect 65313 5200 65335 5400
rect 65486 5200 65513 5400
rect 65514 5200 65541 5400
rect 65692 5200 65714 5400
rect 65720 5200 65742 5400
rect 65893 5200 65920 5400
rect 65921 5200 65948 5400
rect 66099 5200 66121 5400
rect 66127 5200 66149 5400
rect 66300 5200 66327 5400
rect 66328 5200 66355 5400
rect 66506 5200 66528 5400
rect 66534 5200 66556 5400
rect 66707 5200 66734 5400
rect 66735 5200 66762 5400
rect 66913 5200 66935 5400
rect 66941 5200 66963 5400
rect 67114 5200 67141 5400
rect 67142 5200 67169 5400
rect 67320 5200 67342 5400
rect 67348 5200 67370 5400
rect 67521 5200 67548 5400
rect 67549 5200 67576 5400
rect 67727 5200 67749 5400
rect 67755 5200 67777 5400
rect 67928 5200 67955 5400
rect 67956 5200 67983 5400
rect 68134 5200 68156 5400
rect 68162 5200 68184 5400
rect 52869 4800 52896 5000
rect 52897 4800 52924 5000
rect 53070 4800 53097 5000
rect 53098 4800 53125 5000
rect 53271 4800 53298 5000
rect 53299 4800 53326 5000
rect 53477 4800 53499 5000
rect 53505 4800 53527 5000
rect 53683 4800 53705 5000
rect 53711 4800 53733 5000
rect 53884 4800 53911 5000
rect 53912 4800 53939 5000
rect 54085 4800 54112 5000
rect 54113 4800 54140 5000
rect 54291 4800 54313 5000
rect 54319 4800 54341 5000
rect 54497 4800 54519 5000
rect 54525 4800 54547 5000
rect 54703 4800 54725 5000
rect 54731 4800 54753 5000
rect 54904 4800 54931 5000
rect 54932 4800 54959 5000
rect 55110 4800 55132 5000
rect 55138 4800 55160 5000
rect 55311 4800 55338 5000
rect 55339 4800 55366 5000
rect 55517 4800 55539 5000
rect 55545 4800 55567 5000
rect 55718 4800 55745 5000
rect 55746 4800 55773 5000
rect 55924 4800 55946 5000
rect 55952 4800 55974 5000
rect 56125 4800 56152 5000
rect 56153 4800 56180 5000
rect 56331 4800 56353 5000
rect 56359 4800 56381 5000
rect 56532 4800 56559 5000
rect 56560 4800 56587 5000
rect 56738 4800 56760 5000
rect 56766 4800 56788 5000
rect 56944 4800 56966 5000
rect 56972 4800 56994 5000
rect 57145 4800 57172 5000
rect 57173 4800 57200 5000
rect 57346 4800 57373 5000
rect 57374 4800 57401 5000
rect 57552 4800 57574 5000
rect 57580 4800 57602 5000
rect 57753 4800 57780 5000
rect 57781 4800 57808 5000
rect 57959 4800 57981 5000
rect 57987 4800 58009 5000
rect 58160 4800 58187 5000
rect 58188 4800 58215 5000
rect 58366 4800 58388 5000
rect 58394 4800 58416 5000
rect 58567 4800 58594 5000
rect 58595 4800 58622 5000
rect 58773 4800 58795 5000
rect 58801 4800 58823 5000
rect 58974 4800 59001 5000
rect 59002 4800 59029 5000
rect 59180 4800 59202 5000
rect 59208 4800 59230 5000
rect 59381 4800 59408 5000
rect 59409 4800 59436 5000
rect 59587 4800 59609 5000
rect 59615 4800 59637 5000
rect 59788 4800 59815 5000
rect 59816 4800 59843 5000
rect 59994 4800 60016 5000
rect 60022 4800 60044 5000
rect 60195 4800 60222 5000
rect 60223 4800 60250 5000
rect 60401 4800 60423 5000
rect 60429 4800 60451 5000
rect 60602 4800 60629 5000
rect 60630 4800 60657 5000
rect 60808 4800 60830 5000
rect 60836 4800 60858 5000
rect 61009 4800 61036 5000
rect 61037 4800 61064 5000
rect 61215 4800 61237 5000
rect 61243 4800 61265 5000
rect 61416 4800 61443 5000
rect 61444 4800 61471 5000
rect 61622 4800 61644 5000
rect 61650 4800 61672 5000
rect 61823 4800 61850 5000
rect 61851 4800 61878 5000
rect 62029 4800 62051 5000
rect 62057 4800 62079 5000
rect 62230 4800 62257 5000
rect 62258 4800 62285 5000
rect 62436 4800 62458 5000
rect 62464 4800 62486 5000
rect 62637 4800 62664 5000
rect 62665 4800 62692 5000
rect 62843 4800 62865 5000
rect 62871 4800 62893 5000
rect 63044 4800 63071 5000
rect 63072 4800 63099 5000
rect 63250 4800 63272 5000
rect 63278 4800 63300 5000
rect 63451 4800 63478 5000
rect 63479 4800 63506 5000
rect 63657 4800 63679 5000
rect 63685 4800 63707 5000
rect 63858 4800 63885 5000
rect 63886 4800 63913 5000
rect 64064 4800 64086 5000
rect 64092 4800 64114 5000
rect 64265 4800 64292 5000
rect 64293 4800 64320 5000
rect 64471 4800 64493 5000
rect 64499 4800 64521 5000
rect 64672 4800 64699 5000
rect 64700 4800 64727 5000
rect 64878 4800 64900 5000
rect 64906 4800 64928 5000
rect 65079 4800 65106 5000
rect 65107 4800 65134 5000
rect 65285 4800 65307 5000
rect 65313 4800 65335 5000
rect 65486 4800 65513 5000
rect 65514 4800 65541 5000
rect 65692 4800 65714 5000
rect 65720 4800 65742 5000
rect 65893 4800 65920 5000
rect 65921 4800 65948 5000
rect 66099 4800 66121 5000
rect 66127 4800 66149 5000
rect 66300 4800 66327 5000
rect 66328 4800 66355 5000
rect 66506 4800 66528 5000
rect 66534 4800 66556 5000
rect 66707 4800 66734 5000
rect 66735 4800 66762 5000
rect 66913 4800 66935 5000
rect 66941 4800 66963 5000
rect 67114 4800 67141 5000
rect 67142 4800 67169 5000
rect 67320 4800 67342 5000
rect 67348 4800 67370 5000
rect 67521 4800 67548 5000
rect 67549 4800 67576 5000
rect 67727 4800 67749 5000
rect 67755 4800 67777 5000
rect 67928 4800 67955 5000
rect 67956 4800 67983 5000
rect 68134 4800 68156 5000
rect 68162 4800 68184 5000
rect 52869 4400 52896 4600
rect 52897 4400 52924 4600
rect 53070 4400 53097 4600
rect 53098 4400 53125 4600
rect 53271 4400 53298 4600
rect 53299 4400 53326 4600
rect 53477 4400 53499 4600
rect 53505 4400 53527 4600
rect 53683 4400 53705 4600
rect 53711 4400 53733 4600
rect 53884 4400 53911 4600
rect 53912 4400 53939 4600
rect 54085 4400 54112 4600
rect 54113 4400 54140 4600
rect 54291 4400 54313 4600
rect 54319 4400 54341 4600
rect 54497 4400 54519 4600
rect 54525 4400 54547 4600
rect 54703 4400 54725 4600
rect 54731 4400 54753 4600
rect 54904 4400 54931 4600
rect 54932 4400 54959 4600
rect 55110 4400 55132 4600
rect 55138 4400 55160 4600
rect 55311 4400 55338 4600
rect 55339 4400 55366 4600
rect 55517 4400 55539 4600
rect 55545 4400 55567 4600
rect 55718 4400 55745 4600
rect 55746 4400 55773 4600
rect 55924 4400 55946 4600
rect 55952 4400 55974 4600
rect 56125 4400 56152 4600
rect 56153 4400 56180 4600
rect 56331 4400 56353 4600
rect 56359 4400 56381 4600
rect 56532 4400 56559 4600
rect 56560 4400 56587 4600
rect 56738 4400 56760 4600
rect 56766 4400 56788 4600
rect 56944 4400 56966 4600
rect 56972 4400 56994 4600
rect 57145 4400 57172 4600
rect 57173 4400 57200 4600
rect 57346 4400 57373 4600
rect 57374 4400 57401 4600
rect 57552 4400 57574 4600
rect 57580 4400 57602 4600
rect 57753 4400 57780 4600
rect 57781 4400 57808 4600
rect 57959 4400 57981 4600
rect 57987 4400 58009 4600
rect 58160 4400 58187 4600
rect 58188 4400 58215 4600
rect 58366 4400 58388 4600
rect 58394 4400 58416 4600
rect 58567 4400 58594 4600
rect 58595 4400 58622 4600
rect 58773 4400 58795 4600
rect 58801 4400 58823 4600
rect 58974 4400 59001 4600
rect 59002 4400 59029 4600
rect 59180 4400 59202 4600
rect 59208 4400 59230 4600
rect 59381 4400 59408 4600
rect 59409 4400 59436 4600
rect 59587 4400 59609 4600
rect 59615 4400 59637 4600
rect 59788 4400 59815 4600
rect 59816 4400 59843 4600
rect 59994 4400 60016 4600
rect 60022 4400 60044 4600
rect 60195 4400 60222 4600
rect 60223 4400 60250 4600
rect 60401 4400 60423 4600
rect 60429 4400 60451 4600
rect 60602 4400 60629 4600
rect 60630 4400 60657 4600
rect 60808 4400 60830 4600
rect 60836 4400 60858 4600
rect 61009 4400 61036 4600
rect 61037 4400 61064 4600
rect 61215 4400 61237 4600
rect 61243 4400 61265 4600
rect 61416 4400 61443 4600
rect 61444 4400 61471 4600
rect 61622 4400 61644 4600
rect 61650 4400 61672 4600
rect 61823 4400 61850 4600
rect 61851 4400 61878 4600
rect 62029 4400 62051 4600
rect 62057 4400 62079 4600
rect 62230 4400 62257 4600
rect 62258 4400 62285 4600
rect 62436 4400 62458 4600
rect 62464 4400 62486 4600
rect 62637 4400 62664 4600
rect 62665 4400 62692 4600
rect 62843 4400 62865 4600
rect 62871 4400 62893 4600
rect 63044 4400 63071 4600
rect 63072 4400 63099 4600
rect 63250 4400 63272 4600
rect 63278 4400 63300 4600
rect 63451 4400 63478 4600
rect 63479 4400 63506 4600
rect 63657 4400 63679 4600
rect 63685 4400 63707 4600
rect 63858 4400 63885 4600
rect 63886 4400 63913 4600
rect 64064 4400 64086 4600
rect 64092 4400 64114 4600
rect 64265 4400 64292 4600
rect 64293 4400 64320 4600
rect 64471 4400 64493 4600
rect 64499 4400 64521 4600
rect 64672 4400 64699 4600
rect 64700 4400 64727 4600
rect 64878 4400 64900 4600
rect 64906 4400 64928 4600
rect 65079 4400 65106 4600
rect 65107 4400 65134 4600
rect 65285 4400 65307 4600
rect 65313 4400 65335 4600
rect 65486 4400 65513 4600
rect 65514 4400 65541 4600
rect 65692 4400 65714 4600
rect 65720 4400 65742 4600
rect 65893 4400 65920 4600
rect 65921 4400 65948 4600
rect 66099 4400 66121 4600
rect 66127 4400 66149 4600
rect 66300 4400 66327 4600
rect 66328 4400 66355 4600
rect 66506 4400 66528 4600
rect 66534 4400 66556 4600
rect 66707 4400 66734 4600
rect 66735 4400 66762 4600
rect 66913 4400 66935 4600
rect 66941 4400 66963 4600
rect 67114 4400 67141 4600
rect 67142 4400 67169 4600
rect 67320 4400 67342 4600
rect 67348 4400 67370 4600
rect 67521 4400 67548 4600
rect 67549 4400 67576 4600
rect 67727 4400 67749 4600
rect 67755 4400 67777 4600
rect 67928 4400 67955 4600
rect 67956 4400 67983 4600
rect 68134 4400 68156 4600
rect 68162 4400 68184 4600
rect 52869 4000 52896 4200
rect 52897 4000 52924 4200
rect 53070 4000 53097 4200
rect 53098 4000 53125 4200
rect 53271 4000 53298 4200
rect 53299 4000 53326 4200
rect 53477 4000 53499 4200
rect 53505 4000 53527 4200
rect 53683 4000 53705 4200
rect 53711 4000 53733 4200
rect 53884 4000 53911 4200
rect 53912 4000 53939 4200
rect 54085 4000 54112 4200
rect 54113 4000 54140 4200
rect 54291 4000 54313 4200
rect 54319 4000 54341 4200
rect 54497 4000 54519 4200
rect 54525 4000 54547 4200
rect 54703 4000 54725 4200
rect 54731 4000 54753 4200
rect 54904 4000 54931 4200
rect 54932 4000 54959 4200
rect 55110 4000 55132 4200
rect 55138 4000 55160 4200
rect 55311 4000 55338 4200
rect 55339 4000 55366 4200
rect 55517 4000 55539 4200
rect 55545 4000 55567 4200
rect 55718 4000 55745 4200
rect 55746 4000 55773 4200
rect 55924 4000 55946 4200
rect 55952 4000 55974 4200
rect 56125 4000 56152 4200
rect 56153 4000 56180 4200
rect 56331 4000 56353 4200
rect 56359 4000 56381 4200
rect 56532 4000 56559 4200
rect 56560 4000 56587 4200
rect 56738 4000 56760 4200
rect 56766 4000 56788 4200
rect 56944 4000 56966 4200
rect 56972 4000 56994 4200
rect 57145 4000 57172 4200
rect 57173 4000 57200 4200
rect 57346 4000 57373 4200
rect 57374 4000 57401 4200
rect 57552 4000 57574 4200
rect 57580 4000 57602 4200
rect 57753 4000 57780 4200
rect 57781 4000 57808 4200
rect 57959 4000 57981 4200
rect 57987 4000 58009 4200
rect 58160 4000 58187 4200
rect 58188 4000 58215 4200
rect 58366 4000 58388 4200
rect 58394 4000 58416 4200
rect 58567 4000 58594 4200
rect 58595 4000 58622 4200
rect 58773 4000 58795 4200
rect 58801 4000 58823 4200
rect 58974 4000 59001 4200
rect 59002 4000 59029 4200
rect 59180 4000 59202 4200
rect 59208 4000 59230 4200
rect 59381 4000 59408 4200
rect 59409 4000 59436 4200
rect 59587 4000 59609 4200
rect 59615 4000 59637 4200
rect 59788 4000 59815 4200
rect 59816 4000 59843 4200
rect 59994 4000 60016 4200
rect 60022 4000 60044 4200
rect 60195 4000 60222 4200
rect 60223 4000 60250 4200
rect 60401 4000 60423 4200
rect 60429 4000 60451 4200
rect 60602 4000 60629 4200
rect 60630 4000 60657 4200
rect 60808 4000 60830 4200
rect 60836 4000 60858 4200
rect 61009 4000 61036 4200
rect 61037 4000 61064 4200
rect 61215 4000 61237 4200
rect 61243 4000 61265 4200
rect 61416 4000 61443 4200
rect 61444 4000 61471 4200
rect 61622 4000 61644 4200
rect 61650 4000 61672 4200
rect 61823 4000 61850 4200
rect 61851 4000 61878 4200
rect 62029 4000 62051 4200
rect 62057 4000 62079 4200
rect 62230 4000 62257 4200
rect 62258 4000 62285 4200
rect 62436 4000 62458 4200
rect 62464 4000 62486 4200
rect 62637 4000 62664 4200
rect 62665 4000 62692 4200
rect 62843 4000 62865 4200
rect 62871 4000 62893 4200
rect 63044 4000 63071 4200
rect 63072 4000 63099 4200
rect 63250 4000 63272 4200
rect 63278 4000 63300 4200
rect 63451 4000 63478 4200
rect 63479 4000 63506 4200
rect 63657 4000 63679 4200
rect 63685 4000 63707 4200
rect 63858 4000 63885 4200
rect 63886 4000 63913 4200
rect 64064 4000 64086 4200
rect 64092 4000 64114 4200
rect 64265 4000 64292 4200
rect 64293 4000 64320 4200
rect 64471 4000 64493 4200
rect 64499 4000 64521 4200
rect 64672 4000 64699 4200
rect 64700 4000 64727 4200
rect 64878 4000 64900 4200
rect 64906 4000 64928 4200
rect 65079 4000 65106 4200
rect 65107 4000 65134 4200
rect 65285 4000 65307 4200
rect 65313 4000 65335 4200
rect 65486 4000 65513 4200
rect 65514 4000 65541 4200
rect 65692 4000 65714 4200
rect 65720 4000 65742 4200
rect 65893 4000 65920 4200
rect 65921 4000 65948 4200
rect 66099 4000 66121 4200
rect 66127 4000 66149 4200
rect 66300 4000 66327 4200
rect 66328 4000 66355 4200
rect 66506 4000 66528 4200
rect 66534 4000 66556 4200
rect 66707 4000 66734 4200
rect 66735 4000 66762 4200
rect 66913 4000 66935 4200
rect 66941 4000 66963 4200
rect 67114 4000 67141 4200
rect 67142 4000 67169 4200
rect 67320 4000 67342 4200
rect 67348 4000 67370 4200
rect 67521 4000 67548 4200
rect 67549 4000 67576 4200
rect 67727 4000 67749 4200
rect 67755 4000 67777 4200
rect 67928 4000 67955 4200
rect 67956 4000 67983 4200
rect 68134 4000 68156 4200
rect 68162 4000 68184 4200
rect 38382 -1361240 38433 -1361040
rect 38438 -1361240 38461 -1361040
rect 39219 -1361240 39242 -1361040
rect 39247 -1361240 39298 -1361040
rect 39397 -1361240 39448 -1361040
rect 39453 -1361240 39476 -1361040
rect 40033 -1361240 40056 -1361040
rect 40061 -1361240 40112 -1361040
rect 40239 -1361240 40262 -1361040
rect 40267 -1361240 40290 -1361040
rect 40445 -1361240 40468 -1361040
rect 40473 -1361240 40496 -1361040
rect 40852 -1361240 40875 -1361040
rect 40880 -1361240 40903 -1361040
rect 41259 -1361240 41282 -1361040
rect 41287 -1361240 41310 -1361040
rect 41666 -1361240 41689 -1361040
rect 41694 -1361240 41717 -1361040
rect 42073 -1361240 42096 -1361040
rect 42101 -1361240 42124 -1361040
rect 42480 -1361240 42503 -1361040
rect 42508 -1361240 42531 -1361040
rect 42658 -1361240 42709 -1361040
rect 42714 -1361240 42737 -1361040
rect 43294 -1361240 43317 -1361040
rect 43322 -1361240 43373 -1361040
rect 43701 -1361240 43724 -1361040
rect 43729 -1361240 43752 -1361040
rect 44108 -1361240 44131 -1361040
rect 44136 -1361240 44159 -1361040
rect 44515 -1361240 44538 -1361040
rect 44543 -1361240 44566 -1361040
rect 44922 -1361240 44945 -1361040
rect 44950 -1361240 44973 -1361040
rect 45329 -1361240 45352 -1361040
rect 45357 -1361240 45380 -1361040
rect 45736 -1361240 45759 -1361040
rect 45764 -1361240 45787 -1361040
rect 46143 -1361240 46166 -1361040
rect 46171 -1361240 46194 -1361040
rect 46550 -1361240 46573 -1361040
rect 46578 -1361240 46601 -1361040
rect 46957 -1361240 46980 -1361040
rect 46985 -1361240 47008 -1361040
rect 47364 -1361240 47387 -1361040
rect 47392 -1361240 47415 -1361040
rect 47771 -1361240 47794 -1361040
rect 47799 -1361240 47822 -1361040
rect 48178 -1361240 48201 -1361040
rect 48206 -1361240 48229 -1361040
rect 48585 -1361240 48608 -1361040
rect 48613 -1361240 48636 -1361040
rect 48992 -1361240 49015 -1361040
rect 49020 -1361240 49043 -1361040
rect 49399 -1361240 49422 -1361040
rect 49427 -1361240 49450 -1361040
rect 49806 -1361240 49829 -1361040
rect 49834 -1361240 49857 -1361040
rect 50213 -1361240 50236 -1361040
rect 50241 -1361240 50264 -1361040
rect 50620 -1361240 50643 -1361040
rect 50648 -1361240 50671 -1361040
rect 51027 -1361240 51050 -1361040
rect 51055 -1361240 51078 -1361040
rect 51434 -1361240 51457 -1361040
rect 51462 -1361240 51485 -1361040
rect 51841 -1361240 51864 -1361040
rect 51869 -1361240 51892 -1361040
rect 52248 -1361240 52271 -1361040
rect 52276 -1361240 52299 -1361040
rect 52655 -1361240 52678 -1361040
rect 52683 -1361240 52706 -1361040
rect 53062 -1361240 53085 -1361040
rect 53090 -1361240 53113 -1361040
rect 53469 -1361240 53492 -1361040
rect 53497 -1361240 53520 -1361040
rect 53876 -1361240 53899 -1361040
rect 53904 -1361240 53927 -1361040
rect 38382 -1361640 38433 -1361440
rect 38438 -1361640 38461 -1361440
rect 39219 -1361640 39242 -1361440
rect 39247 -1361640 39298 -1361440
rect 39397 -1361640 39448 -1361440
rect 39453 -1361640 39476 -1361440
rect 40033 -1361640 40056 -1361440
rect 40061 -1361640 40112 -1361440
rect 40239 -1361640 40262 -1361440
rect 40267 -1361640 40290 -1361440
rect 40445 -1361640 40468 -1361440
rect 40473 -1361640 40496 -1361440
rect 40852 -1361640 40875 -1361440
rect 40880 -1361640 40903 -1361440
rect 41259 -1361640 41282 -1361440
rect 41287 -1361640 41310 -1361440
rect 41666 -1361640 41689 -1361440
rect 41694 -1361640 41717 -1361440
rect 42073 -1361640 42096 -1361440
rect 42101 -1361640 42124 -1361440
rect 42480 -1361640 42503 -1361440
rect 42508 -1361640 42531 -1361440
rect 42658 -1361640 42709 -1361440
rect 42714 -1361640 42737 -1361440
rect 43294 -1361640 43317 -1361440
rect 43322 -1361640 43373 -1361440
rect 43701 -1361640 43724 -1361440
rect 43729 -1361640 43752 -1361440
rect 44108 -1361640 44131 -1361440
rect 44136 -1361640 44159 -1361440
rect 44515 -1361640 44538 -1361440
rect 44543 -1361640 44566 -1361440
rect 44922 -1361640 44945 -1361440
rect 44950 -1361640 44973 -1361440
rect 45329 -1361640 45352 -1361440
rect 45357 -1361640 45380 -1361440
rect 45736 -1361640 45759 -1361440
rect 45764 -1361640 45787 -1361440
rect 46143 -1361640 46166 -1361440
rect 46171 -1361640 46194 -1361440
rect 46550 -1361640 46573 -1361440
rect 46578 -1361640 46601 -1361440
rect 46957 -1361640 46980 -1361440
rect 46985 -1361640 47008 -1361440
rect 47364 -1361640 47387 -1361440
rect 47392 -1361640 47415 -1361440
rect 47771 -1361640 47794 -1361440
rect 47799 -1361640 47822 -1361440
rect 48178 -1361640 48201 -1361440
rect 48206 -1361640 48229 -1361440
rect 48585 -1361640 48608 -1361440
rect 48613 -1361640 48636 -1361440
rect 48992 -1361640 49015 -1361440
rect 49020 -1361640 49043 -1361440
rect 49399 -1361640 49422 -1361440
rect 49427 -1361640 49450 -1361440
rect 49806 -1361640 49829 -1361440
rect 49834 -1361640 49857 -1361440
rect 50213 -1361640 50236 -1361440
rect 50241 -1361640 50264 -1361440
rect 50620 -1361640 50643 -1361440
rect 50648 -1361640 50671 -1361440
rect 51027 -1361640 51050 -1361440
rect 51055 -1361640 51078 -1361440
rect 51434 -1361640 51457 -1361440
rect 51462 -1361640 51485 -1361440
rect 51841 -1361640 51864 -1361440
rect 51869 -1361640 51892 -1361440
rect 52248 -1361640 52271 -1361440
rect 52276 -1361640 52299 -1361440
rect 52655 -1361640 52678 -1361440
rect 52683 -1361640 52706 -1361440
rect 53062 -1361640 53085 -1361440
rect 53090 -1361640 53113 -1361440
rect 53469 -1361640 53492 -1361440
rect 53497 -1361640 53520 -1361440
rect 53876 -1361640 53899 -1361440
rect 53904 -1361640 53927 -1361440
rect 38382 -1362040 38433 -1361840
rect 38438 -1362040 38461 -1361840
rect 39219 -1362040 39242 -1361840
rect 39247 -1362040 39298 -1361840
rect 39397 -1362040 39448 -1361840
rect 39453 -1362040 39476 -1361840
rect 40033 -1362040 40056 -1361840
rect 40061 -1362040 40112 -1361840
rect 40239 -1362040 40262 -1361840
rect 40267 -1362040 40290 -1361840
rect 40445 -1362040 40468 -1361840
rect 40473 -1362040 40496 -1361840
rect 40852 -1362040 40875 -1361840
rect 40880 -1362040 40903 -1361840
rect 41259 -1362040 41282 -1361840
rect 41287 -1362040 41310 -1361840
rect 41666 -1362040 41689 -1361840
rect 41694 -1362040 41717 -1361840
rect 42073 -1362040 42096 -1361840
rect 42101 -1362040 42124 -1361840
rect 42480 -1362040 42503 -1361840
rect 42508 -1362040 42531 -1361840
rect 42658 -1362040 42709 -1361840
rect 42714 -1362040 42737 -1361840
rect 43294 -1362040 43317 -1361840
rect 43322 -1362040 43373 -1361840
rect 43701 -1362040 43724 -1361840
rect 43729 -1362040 43752 -1361840
rect 44108 -1362040 44131 -1361840
rect 44136 -1362040 44159 -1361840
rect 44515 -1362040 44538 -1361840
rect 44543 -1362040 44566 -1361840
rect 44922 -1362040 44945 -1361840
rect 44950 -1362040 44973 -1361840
rect 45329 -1362040 45352 -1361840
rect 45357 -1362040 45380 -1361840
rect 45736 -1362040 45759 -1361840
rect 45764 -1362040 45787 -1361840
rect 46143 -1362040 46166 -1361840
rect 46171 -1362040 46194 -1361840
rect 46550 -1362040 46573 -1361840
rect 46578 -1362040 46601 -1361840
rect 46957 -1362040 46980 -1361840
rect 46985 -1362040 47008 -1361840
rect 47364 -1362040 47387 -1361840
rect 47392 -1362040 47415 -1361840
rect 47771 -1362040 47794 -1361840
rect 47799 -1362040 47822 -1361840
rect 48178 -1362040 48201 -1361840
rect 48206 -1362040 48229 -1361840
rect 48585 -1362040 48608 -1361840
rect 48613 -1362040 48636 -1361840
rect 48992 -1362040 49015 -1361840
rect 49020 -1362040 49043 -1361840
rect 49399 -1362040 49422 -1361840
rect 49427 -1362040 49450 -1361840
rect 49806 -1362040 49829 -1361840
rect 49834 -1362040 49857 -1361840
rect 50213 -1362040 50236 -1361840
rect 50241 -1362040 50264 -1361840
rect 50620 -1362040 50643 -1361840
rect 50648 -1362040 50671 -1361840
rect 51027 -1362040 51050 -1361840
rect 51055 -1362040 51078 -1361840
rect 51434 -1362040 51457 -1361840
rect 51462 -1362040 51485 -1361840
rect 51841 -1362040 51864 -1361840
rect 51869 -1362040 51892 -1361840
rect 52248 -1362040 52271 -1361840
rect 52276 -1362040 52299 -1361840
rect 52655 -1362040 52678 -1361840
rect 52683 -1362040 52706 -1361840
rect 53062 -1362040 53085 -1361840
rect 53090 -1362040 53113 -1361840
rect 53469 -1362040 53492 -1361840
rect 53497 -1362040 53520 -1361840
rect 53876 -1362040 53899 -1361840
rect 53904 -1362040 53927 -1361840
rect 39219 -1362440 39242 -1362240
rect 39247 -1362440 39298 -1362240
rect 39397 -1362440 39448 -1362240
rect 39453 -1362440 39476 -1362240
rect 40033 -1362440 40056 -1362240
rect 40061 -1362440 40112 -1362240
rect 40239 -1362440 40262 -1362240
rect 40267 -1362440 40290 -1362240
rect 40445 -1362440 40468 -1362240
rect 40473 -1362440 40496 -1362240
rect 40852 -1362440 40875 -1362240
rect 40880 -1362440 40903 -1362240
rect 41259 -1362440 41282 -1362240
rect 41287 -1362440 41310 -1362240
rect 41666 -1362440 41689 -1362240
rect 41694 -1362440 41717 -1362240
rect 42073 -1362440 42096 -1362240
rect 42101 -1362440 42124 -1362240
rect 42480 -1362440 42503 -1362240
rect 42508 -1362440 42531 -1362240
rect 42658 -1362440 42709 -1362240
rect 42714 -1362440 42737 -1362240
rect 43294 -1362440 43317 -1362240
rect 43322 -1362440 43373 -1362240
rect 43701 -1362440 43724 -1362240
rect 43729 -1362440 43752 -1362240
rect 44108 -1362440 44131 -1362240
rect 44136 -1362440 44159 -1362240
rect 44515 -1362440 44538 -1362240
rect 44543 -1362440 44566 -1362240
rect 44922 -1362440 44945 -1362240
rect 44950 -1362440 44973 -1362240
rect 45329 -1362440 45352 -1362240
rect 45357 -1362440 45380 -1362240
rect 45736 -1362440 45759 -1362240
rect 45764 -1362440 45787 -1362240
rect 46143 -1362440 46166 -1362240
rect 46171 -1362440 46194 -1362240
rect 46550 -1362440 46573 -1362240
rect 46578 -1362440 46601 -1362240
rect 46957 -1362440 46980 -1362240
rect 46985 -1362440 47008 -1362240
rect 47364 -1362440 47387 -1362240
rect 47392 -1362440 47415 -1362240
rect 47771 -1362440 47794 -1362240
rect 47799 -1362440 47822 -1362240
rect 48178 -1362440 48201 -1362240
rect 48206 -1362440 48229 -1362240
rect 48585 -1362440 48608 -1362240
rect 48613 -1362440 48636 -1362240
rect 48992 -1362440 49015 -1362240
rect 49020 -1362440 49043 -1362240
rect 49399 -1362440 49422 -1362240
rect 49427 -1362440 49450 -1362240
rect 49806 -1362440 49829 -1362240
rect 49834 -1362440 49857 -1362240
rect 50213 -1362440 50236 -1362240
rect 50241 -1362440 50264 -1362240
rect 50620 -1362440 50643 -1362240
rect 50648 -1362440 50671 -1362240
rect 51027 -1362440 51050 -1362240
rect 51055 -1362440 51078 -1362240
rect 51434 -1362440 51457 -1362240
rect 51462 -1362440 51485 -1362240
rect 51841 -1362440 51864 -1362240
rect 51869 -1362440 51892 -1362240
rect 52248 -1362440 52271 -1362240
rect 52276 -1362440 52299 -1362240
rect 52655 -1362440 52678 -1362240
rect 52683 -1362440 52706 -1362240
rect 53062 -1362440 53085 -1362240
rect 53090 -1362440 53113 -1362240
rect 53469 -1362440 53492 -1362240
rect 53497 -1362440 53520 -1362240
rect 53876 -1362440 53899 -1362240
rect 53904 -1362440 53927 -1362240
rect 39219 -1362840 39242 -1362640
rect 39247 -1362840 39298 -1362640
rect 39397 -1362840 39448 -1362640
rect 39453 -1362840 39476 -1362640
rect 40033 -1362840 40056 -1362640
rect 40061 -1362840 40112 -1362640
rect 40239 -1362840 40262 -1362640
rect 40267 -1362840 40290 -1362640
rect 40445 -1362840 40468 -1362640
rect 40473 -1362840 40496 -1362640
rect 40852 -1362840 40875 -1362640
rect 40880 -1362840 40903 -1362640
rect 41259 -1362840 41282 -1362640
rect 41287 -1362840 41310 -1362640
rect 41666 -1362840 41689 -1362640
rect 41694 -1362840 41717 -1362640
rect 42073 -1362840 42096 -1362640
rect 42101 -1362840 42124 -1362640
rect 42480 -1362840 42503 -1362640
rect 42508 -1362840 42531 -1362640
rect 42658 -1362840 42709 -1362640
rect 42714 -1362840 42737 -1362640
rect 43294 -1362840 43317 -1362640
rect 43322 -1362840 43373 -1362640
rect 43701 -1362840 43724 -1362640
rect 43729 -1362840 43752 -1362640
rect 44108 -1362840 44131 -1362640
rect 44136 -1362840 44159 -1362640
rect 44515 -1362840 44538 -1362640
rect 44543 -1362840 44566 -1362640
rect 44922 -1362840 44945 -1362640
rect 44950 -1362840 44973 -1362640
rect 45329 -1362840 45352 -1362640
rect 45357 -1362840 45380 -1362640
rect 45736 -1362840 45759 -1362640
rect 45764 -1362840 45787 -1362640
rect 46143 -1362840 46166 -1362640
rect 46171 -1362840 46194 -1362640
rect 46550 -1362840 46573 -1362640
rect 46578 -1362840 46601 -1362640
rect 46957 -1362840 46980 -1362640
rect 46985 -1362840 47008 -1362640
rect 47364 -1362840 47387 -1362640
rect 47392 -1362840 47415 -1362640
rect 47771 -1362840 47794 -1362640
rect 47799 -1362840 47822 -1362640
rect 48178 -1362840 48201 -1362640
rect 48206 -1362840 48229 -1362640
rect 48585 -1362840 48608 -1362640
rect 48613 -1362840 48636 -1362640
rect 48992 -1362840 49015 -1362640
rect 49020 -1362840 49043 -1362640
rect 49399 -1362840 49422 -1362640
rect 49427 -1362840 49450 -1362640
rect 49806 -1362840 49829 -1362640
rect 49834 -1362840 49857 -1362640
rect 50213 -1362840 50236 -1362640
rect 50241 -1362840 50264 -1362640
rect 50620 -1362840 50643 -1362640
rect 50648 -1362840 50671 -1362640
rect 51027 -1362840 51050 -1362640
rect 51055 -1362840 51078 -1362640
rect 51434 -1362840 51457 -1362640
rect 51462 -1362840 51485 -1362640
rect 51841 -1362840 51864 -1362640
rect 51869 -1362840 51892 -1362640
rect 52248 -1362840 52271 -1362640
rect 52276 -1362840 52299 -1362640
rect 52655 -1362840 52678 -1362640
rect 52683 -1362840 52706 -1362640
rect 53062 -1362840 53085 -1362640
rect 53090 -1362840 53113 -1362640
rect 53469 -1362840 53492 -1362640
rect 53497 -1362840 53520 -1362640
rect 53876 -1362840 53899 -1362640
rect 53904 -1362840 53927 -1362640
rect 39219 -1363240 39242 -1363040
rect 39247 -1363240 39298 -1363040
rect 39397 -1363240 39448 -1363040
rect 39453 -1363240 39476 -1363040
rect 40033 -1363240 40056 -1363040
rect 40061 -1363240 40112 -1363040
rect 40239 -1363240 40262 -1363040
rect 40267 -1363240 40290 -1363040
rect 40445 -1363240 40468 -1363040
rect 40473 -1363240 40496 -1363040
rect 40852 -1363240 40875 -1363040
rect 40880 -1363240 40903 -1363040
rect 41259 -1363240 41282 -1363040
rect 41287 -1363240 41310 -1363040
rect 41666 -1363240 41689 -1363040
rect 41694 -1363240 41717 -1363040
rect 42073 -1363240 42096 -1363040
rect 42101 -1363240 42124 -1363040
rect 42480 -1363240 42503 -1363040
rect 42508 -1363240 42531 -1363040
rect 42658 -1363240 42709 -1363040
rect 42714 -1363240 42737 -1363040
rect 43294 -1363240 43317 -1363040
rect 43322 -1363240 43373 -1363040
rect 43701 -1363240 43724 -1363040
rect 43729 -1363240 43752 -1363040
rect 44108 -1363240 44131 -1363040
rect 44136 -1363240 44159 -1363040
rect 44515 -1363240 44538 -1363040
rect 44543 -1363240 44566 -1363040
rect 44922 -1363240 44945 -1363040
rect 44950 -1363240 44973 -1363040
rect 45329 -1363240 45352 -1363040
rect 45357 -1363240 45380 -1363040
rect 45736 -1363240 45759 -1363040
rect 45764 -1363240 45787 -1363040
rect 46143 -1363240 46166 -1363040
rect 46171 -1363240 46194 -1363040
rect 46550 -1363240 46573 -1363040
rect 46578 -1363240 46601 -1363040
rect 46957 -1363240 46980 -1363040
rect 46985 -1363240 47008 -1363040
rect 47364 -1363240 47387 -1363040
rect 47392 -1363240 47415 -1363040
rect 47771 -1363240 47794 -1363040
rect 47799 -1363240 47822 -1363040
rect 48178 -1363240 48201 -1363040
rect 48206 -1363240 48229 -1363040
rect 48585 -1363240 48608 -1363040
rect 48613 -1363240 48636 -1363040
rect 48992 -1363240 49015 -1363040
rect 49020 -1363240 49043 -1363040
rect 49399 -1363240 49422 -1363040
rect 49427 -1363240 49450 -1363040
rect 49806 -1363240 49829 -1363040
rect 49834 -1363240 49857 -1363040
rect 50213 -1363240 50236 -1363040
rect 50241 -1363240 50264 -1363040
rect 50620 -1363240 50643 -1363040
rect 50648 -1363240 50671 -1363040
rect 51027 -1363240 51050 -1363040
rect 51055 -1363240 51078 -1363040
rect 51434 -1363240 51457 -1363040
rect 51462 -1363240 51485 -1363040
rect 51841 -1363240 51864 -1363040
rect 51869 -1363240 51892 -1363040
rect 52248 -1363240 52271 -1363040
rect 52276 -1363240 52299 -1363040
rect 52655 -1363240 52678 -1363040
rect 52683 -1363240 52706 -1363040
rect 53062 -1363240 53085 -1363040
rect 53090 -1363240 53113 -1363040
rect 53469 -1363240 53492 -1363040
rect 53497 -1363240 53520 -1363040
rect 53876 -1363240 53899 -1363040
rect 53904 -1363240 53927 -1363040
rect 39219 -1363640 39242 -1363440
rect 39247 -1363640 39298 -1363440
rect 39397 -1363640 39448 -1363440
rect 39453 -1363640 39476 -1363440
rect 40033 -1363640 40056 -1363440
rect 40061 -1363640 40112 -1363440
rect 40239 -1363640 40262 -1363440
rect 40267 -1363640 40290 -1363440
rect 40445 -1363640 40468 -1363440
rect 40473 -1363640 40496 -1363440
rect 40852 -1363640 40875 -1363440
rect 40880 -1363640 40903 -1363440
rect 41259 -1363640 41282 -1363440
rect 41287 -1363640 41310 -1363440
rect 41666 -1363640 41689 -1363440
rect 41694 -1363640 41717 -1363440
rect 42073 -1363640 42096 -1363440
rect 42101 -1363640 42124 -1363440
rect 42480 -1363640 42503 -1363440
rect 42508 -1363640 42531 -1363440
rect 42658 -1363640 42709 -1363440
rect 42714 -1363640 42737 -1363440
rect 43294 -1363640 43317 -1363440
rect 43322 -1363640 43373 -1363440
rect 43701 -1363640 43724 -1363440
rect 43729 -1363640 43752 -1363440
rect 44108 -1363640 44131 -1363440
rect 44136 -1363640 44159 -1363440
rect 44515 -1363640 44538 -1363440
rect 44543 -1363640 44566 -1363440
rect 44922 -1363640 44945 -1363440
rect 44950 -1363640 44973 -1363440
rect 45329 -1363640 45352 -1363440
rect 45357 -1363640 45380 -1363440
rect 45736 -1363640 45759 -1363440
rect 45764 -1363640 45787 -1363440
rect 46143 -1363640 46166 -1363440
rect 46171 -1363640 46194 -1363440
rect 46550 -1363640 46573 -1363440
rect 46578 -1363640 46601 -1363440
rect 46957 -1363640 46980 -1363440
rect 46985 -1363640 47008 -1363440
rect 47364 -1363640 47387 -1363440
rect 47392 -1363640 47415 -1363440
rect 47771 -1363640 47794 -1363440
rect 47799 -1363640 47822 -1363440
rect 48178 -1363640 48201 -1363440
rect 48206 -1363640 48229 -1363440
rect 48585 -1363640 48608 -1363440
rect 48613 -1363640 48636 -1363440
rect 48992 -1363640 49015 -1363440
rect 49020 -1363640 49043 -1363440
rect 49399 -1363640 49422 -1363440
rect 49427 -1363640 49450 -1363440
rect 49806 -1363640 49829 -1363440
rect 49834 -1363640 49857 -1363440
rect 50213 -1363640 50236 -1363440
rect 50241 -1363640 50264 -1363440
rect 50620 -1363640 50643 -1363440
rect 50648 -1363640 50671 -1363440
rect 51027 -1363640 51050 -1363440
rect 51055 -1363640 51078 -1363440
rect 51434 -1363640 51457 -1363440
rect 51462 -1363640 51485 -1363440
rect 51841 -1363640 51864 -1363440
rect 51869 -1363640 51892 -1363440
rect 52248 -1363640 52271 -1363440
rect 52276 -1363640 52299 -1363440
rect 52655 -1363640 52678 -1363440
rect 52683 -1363640 52706 -1363440
rect 53062 -1363640 53085 -1363440
rect 53090 -1363640 53113 -1363440
rect 53469 -1363640 53492 -1363440
rect 53497 -1363640 53520 -1363440
rect 53876 -1363640 53899 -1363440
rect 53904 -1363640 53927 -1363440
rect 39219 -1364040 39242 -1363840
rect 39247 -1364040 39270 -1363840
rect 39425 -1364040 39448 -1363840
rect 39453 -1364040 39476 -1363840
rect 40033 -1364040 40056 -1363840
rect 40061 -1364040 40084 -1363840
rect 40239 -1364040 40262 -1363840
rect 40267 -1364040 40290 -1363840
rect 40445 -1364040 40468 -1363840
rect 40473 -1364040 40496 -1363840
rect 40852 -1364040 40875 -1363840
rect 40880 -1364040 40903 -1363840
rect 41259 -1364040 41282 -1363840
rect 41287 -1364040 41310 -1363840
rect 41666 -1364040 41689 -1363840
rect 41694 -1364040 41717 -1363840
rect 42073 -1364040 42096 -1363840
rect 42101 -1364040 42124 -1363840
rect 42480 -1364040 42503 -1363840
rect 42508 -1364040 42531 -1363840
rect 42686 -1364040 42709 -1363840
rect 42714 -1364040 42737 -1363840
rect 43294 -1364040 43317 -1363840
rect 43322 -1364040 43345 -1363840
rect 43701 -1364040 43724 -1363840
rect 43729 -1364040 43752 -1363840
rect 44108 -1364040 44131 -1363840
rect 44136 -1364040 44159 -1363840
rect 44515 -1364040 44538 -1363840
rect 44543 -1364040 44566 -1363840
rect 44922 -1364040 44945 -1363840
rect 44950 -1364040 44973 -1363840
rect 45329 -1364040 45352 -1363840
rect 45357 -1364040 45380 -1363840
rect 45736 -1364040 45759 -1363840
rect 45764 -1364040 45787 -1363840
rect 46143 -1364040 46166 -1363840
rect 46171 -1364040 46194 -1363840
rect 46550 -1364040 46573 -1363840
rect 46578 -1364040 46601 -1363840
rect 46957 -1364040 46980 -1363840
rect 46985 -1364040 47008 -1363840
rect 47364 -1364040 47387 -1363840
rect 47392 -1364040 47415 -1363840
rect 47771 -1364040 47794 -1363840
rect 47799 -1364040 47822 -1363840
rect 48178 -1364040 48201 -1363840
rect 48206 -1364040 48229 -1363840
rect 48585 -1364040 48608 -1363840
rect 48613 -1364040 48636 -1363840
rect 48992 -1364040 49015 -1363840
rect 49020 -1364040 49043 -1363840
rect 49399 -1364040 49422 -1363840
rect 49427 -1364040 49450 -1363840
rect 49806 -1364040 49829 -1363840
rect 49834 -1364040 49857 -1363840
rect 50213 -1364040 50236 -1363840
rect 50241 -1364040 50264 -1363840
rect 50620 -1364040 50643 -1363840
rect 50648 -1364040 50671 -1363840
rect 51027 -1364040 51050 -1363840
rect 51055 -1364040 51078 -1363840
rect 51434 -1364040 51457 -1363840
rect 51462 -1364040 51485 -1363840
rect 51841 -1364040 51864 -1363840
rect 51869 -1364040 51892 -1363840
rect 52248 -1364040 52271 -1363840
rect 52276 -1364040 52299 -1363840
rect 52655 -1364040 52678 -1363840
rect 52683 -1364040 52706 -1363840
rect 53062 -1364040 53085 -1363840
rect 53090 -1364040 53113 -1363840
rect 53469 -1364040 53492 -1363840
rect 53497 -1364040 53520 -1363840
rect 53876 -1364040 53899 -1363840
rect 53904 -1364040 53927 -1363840
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
use CNR_GR06  CNR_GR06_0
timestamp 1713381030
transform 1 0 0 0 1 2600
box 0 -2000 17197 5531
use CNR_GR06_I_to_t  CNR_GR06_I_to_t_0
timestamp 1713381165
transform 1 0 14258 0 1 1368640
box 0 -1368204 55098 200
use CNR_GR06_I_to_t  CNR_GR06_I_to_t_1
timestamp 1713381165
transform 1 0 0 0 1 600
box 0 -1368204 55098 200
use comparator  comparator_0
timestamp 1713380703
transform 1 0 62681 0 1 3000
box 0 -2400 7251 2767
use comparator  comparator_1
timestamp 1713380703
transform 1 0 58037 0 1 -1365040
box 0 -2400 7251 2767
use comparator  comparator_2
timestamp 1713380703
transform 1 0 2939 0 1 -1365204
box 0 -2400 7251 2767
use dac  dac_0
timestamp 1713380703
transform 1 0 59742 0 1 2200
box 0 -1600 2939 2767
use dac  dac_1
timestamp 1713380703
transform 1 0 55098 0 1 -1365840
box 0 -1600 2939 2767
use dac  dac_2
timestamp 1713380703
transform 1 0 0 0 1 -1366004
box 0 -1600 2939 2767
use dac_n  dac_n_0
timestamp 1713380703
transform 1 0 69932 0 1 2200
box 0 -1600 2939 2767
use dac_n  dac_n_1
timestamp 1713380703
transform 1 0 65288 0 1 -1365840
box 0 -1600 2939 2767
use dac_n  dac_n_2
timestamp 1713380703
transform 1 0 10190 0 1 -1366004
box 0 -1600 2939 2767
use CNR_GR06  x1
timestamp 1713381030
transform 1 0 0 0 1 600
box 0 -2000 17197 5531
use CNR_GR06_I_to_t  x2
timestamp 1713381165
transform 1 0 1 0 1 600
box 0 -1368204 55098 200
use comparator  x3
timestamp 1713380703
transform 1 0 3 0 1 600
box 0 -2400 7251 2767
use dac_n  x4
timestamp 1713380703
transform 1 0 4 0 1 600
box 0 -1600 2939 2767
use dac  x5
timestamp 1713380703
transform 1 0 2 0 1 600
box 0 -1600 2939 2767
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD_1V8
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vn
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vp
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 Vop
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Von
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Clk_1
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 Clk_2
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 Clk
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 VT1
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 VT2
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 Vocn
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 DACN
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 DACP
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 Vdref
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 VBN
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 {}
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 VBP
port 17 nsew
<< end >>
