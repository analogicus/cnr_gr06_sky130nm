* This is your template.sp file

* Other SPICE commands...

.param vth0_n = 
.param vth0_p = 

* More SPICE commands...

